library IEEE;
use IEEE.std_logic_1164.all;  -- defines std_logic types
use IEEE.STD_LOGIC_unsigned.all;
use IEEE.STD_LOGIC_arith.all;

-- microcode 65C816
-- Written by Valerio Venturi
-- output fields format:
-- fields:
-- RSEL:  registers output multiplexer select
-- REGOP: registers load/increment/decrement etc.
-- ALUOP: ALU operation
-- P_OP:  register P set/reset bit
-- MPR:   register MP 
-- PCR:   register PC 
-- CLI:   clear interrupt request
-- EI:    end of microcode sequence
-- W:     read/write control
-- PD:    PC/MP output multiplexer select
-- VPA:   valid program address
-- VDA:   valid data address
-- ML:    memory lock
entity mcpla is
  port(em:  in STD_LOGIC;                           -- emulation mode (1)/native mode (0)
        m:  in STD_LOGIC;                           -- M memory/acc. 8 bit (1), M memory/acc. 16 bit (0)  
        x:  in STD_LOGIC;                           -- X index reg. 8 bit (1), X index reg. 16 bit (0)  
        a:  in STD_LOGIC_VECTOR(12 downto 0);
        q: out STD_LOGIC_VECTOR(44 downto 0)
      );
end mcpla;

architecture comb of mcpla is

constant  MC_ADDR_LENGTH: INTEGER := 12; 
-- opcode definition:
-- <EXPANSION OPCODE (1 BIT) (WDM)>-<OPCODE (8 bits)>-<MICROCODE (4 BITS)>

------------------------------------
--            IMPLIED             --
------------------------------------
constant   NOP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111010100000"; -- 0xEA NOP

-- interrupts/coprocessor
constant   BRK_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000000"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000001"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000010"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000011"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000100"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000101"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000110"; -- 0x00 BRK/IRQ/NMI/RES
constant   BRK_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000000111"; -- 0x00 BRK/IRQ/NMI/RES

constant   COP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100000"; -- 0x02 COP
constant   COP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100001"; -- 0x02 COP
constant   COP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100010"; -- 0x02 COP
constant   COP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100011"; -- 0x02 COP
constant   COP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100100"; -- 0x02 COP
constant   COP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100101"; -- 0x02 COP
constant   COP_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100110"; -- 0x02 COP
constant   COP_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000100111"; -- 0x02 COP

-- IMPLIED
constant   CLC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110000000"; -- 0x18 CLC 0->C 
constant   SEC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110000000"; -- 0x38 SEC 1->C
constant   CLI_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110000000"; -- 0x58 CLI 0->I
constant   SEI_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110000000"; -- 0x78 SEI 1->I
constant   CLV_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110000000"; -- 0xB8 CLV 0->V
constant   CLD_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110000000"; -- 0xD8 CLD 0->D
constant   SED_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110000000"; -- 0xF8 SED 1->D
constant   TAX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101010100000"; -- 0xAA TAX A->X
constant   TAY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101010000000"; -- 0xA8 TAY A->Y
constant   TXA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010100000"; -- 0x8A TXA X->A
constant   TYA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110000000"; -- 0x98 TYA Y->A
constant   TXY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110110000"; -- 0x9B TXY X->Y
constant   TYX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110110000"; -- 0xBB TYX Y->X
constant   TXS_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110100000"; -- 0x9A TXS X->S
constant   TSX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110100000"; -- 0xBA TSX S->X
constant   TCD_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110110000"; -- 0x5B TCD C->D
constant   TDC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110110000"; -- 0x7B TDC D->C
constant   PHP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000010000000"; -- 0x08 PHP P->S
constant   PHA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010010000000"; -- 0x48 PHA A->S
constant   PHA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010010000001"; -- 0x48 PHA A->S
constant   PHX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110100000"; -- 0xDA PHX X->S
constant   PHX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110100001"; -- 0xDA PHX X->S
constant   PHY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110100000"; -- 0x5A PHY X->S
constant   PHY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110100001"; -- 0x5A PHY X->S
constant   PHD_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000010110000"; -- 0x0B PHD D->S
constant   PHD_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000010110001"; -- 0x0B PHD D->S
constant   PLP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010000000"; -- 0x28 PLP S->P
constant   PLP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010000001"; -- 0x28 PLP S->P
constant   PLA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010000000"; -- 0x68 PLA S->A
constant   PLA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010000001"; -- 0x68 PLA S->A
constant   PLA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010000010"; -- 0x68 PLA S->A
constant   PLA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010000011"; -- 0x68 PLA S->A
constant   PLX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110100000"; -- 0xFA PLX S->X
constant   PLX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110100001"; -- 0xFA PLX S->X
constant   PLX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110100010"; -- 0xFA PLX S->X
constant   PLX_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110100011"; -- 0xFA PLX S->X
constant   PLY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110100000"; -- 0x7A PLY S->Y
constant   PLY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110100001"; -- 0x7A PLY S->Y
constant   PLY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110100010"; -- 0x7A PLY S->Y
constant   PLY_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110100011"; -- 0x7A PLY S->Y
constant   PLD_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010110000"; -- 0x2B PLD S->D
constant   PLD_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010110001"; -- 0x2B PLD S->D
constant   PLD_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010110010"; -- 0x2B PLD S->D
constant   INC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110100000"; -- 0x1A INC A +1
constant   DEC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110100000"; -- 0x3A DEC A -1
constant   INX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111010000000"; -- 0xE8 INX X +1
constant   DEX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110010100000"; -- 0xCA DEX X -1
constant   INY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110010000000"; -- 0xC8 INY Y +1
constant   DEY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010000000"; -- 0x88 DEY Y -1
constant   RTS_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000000000"; -- 0x60 RTS    
constant   RTS_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000000001"; -- 0x60 RTS    
constant   RTS_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000000010"; -- 0x60 RTS    
constant   RTS_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000000011"; -- 0x60 RTS    
constant   RTS_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000000100"; -- 0x60 RTS    
constant   RTI_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000000"; -- 0x40 RTI    
constant   RTI_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000001"; -- 0x40 RTI    
constant   RTI_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000010"; -- 0x40 RTI    
constant   RTI_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000011"; -- 0x40 RTI    
constant   RTI_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000100"; -- 0x40 RTI    
constant   RTI_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000101"; -- 0x40 RTI    
constant   RTI_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000000110"; -- 0x40 RTI    
constant   ASL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000010100000"; -- 0x0A ASL A  
constant   LSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010010100000"; -- 0x4A LSR A  
constant   ROL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010100000"; -- 0x2A ROL A  
constant   ROR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010100000"; -- 0x6A ROR A  
constant   TCS_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110110000"; -- 0x1B A->S
constant   TSC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110110000"; -- 0x3B S->A
constant   XCE_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110110000"; -- 0xFB XCE E<->C 
constant   WDM_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000100000"; -- 0x42 WDM
constant   PHK_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010010110000"; -- 0x4B PHK K->S
constant   PHB_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010110000"; -- 0x8B PHB B->S
constant   PLB_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101010110000"; -- 0xAB PLB S->B
constant   PLB_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101010110001"; -- 0xAB PLB S->B
constant   RTL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110000"; -- 0x6B RTL    
constant   RTL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110001"; -- 0x6B RTL    
constant   RTL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110010"; -- 0x6B RTL    
constant   RTL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110011"; -- 0x6B RTL    
constant   RTL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110100"; -- 0x6B RTL    
constant   RTL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110101"; -- 0x6B RTL    
constant   RTL_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010110110"; -- 0x6B RTL    
constant   XBA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111010110000"; -- 0xEB XBA (swap A)
constant   WAI_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110010110000"; -- 0xCB WAI
constant   WAI_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110010110001"; -- 0xCB WAI
constant   STP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110110000"; -- 0xDB STP
constant   STP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110110001"; -- 0xDB STP

------------------------------------
--           IMMEDIATE            --
------------------------------------
constant IMLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101010010000"; -- 0xA9 LDA #IMM
constant IMLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101010010001"; -- 0xA9 LDA #IMM
constant IMLDX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000100000"; -- 0xA2 LDX #IMM
constant IMLDX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000100001"; -- 0xA2 LDX #IMM
constant IMLDY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000000000"; -- 0xA0 LDY #IMM
constant IMLDY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000000001"; -- 0xA0 LDY #IMM
constant IMADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010010000"; -- 0x69 ADC #IMM 
constant IMADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010010001"; -- 0x69 ADC #IMM 
constant IMADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011010010010"; -- 0x69 ADC #IMM 
constant IMSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111010010000"; -- 0xE9 SBC #IMM 
constant IMSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111010010001"; -- 0xE9 SBC #IMM 
constant IMSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111010010010"; -- 0xE9 SBC #IMM 
constant IMAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010010000"; -- 0x29 AND #IMM 
constant IMAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001010010001"; -- 0x29 AND #IMM 
constant IMORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000010010000"; -- 0x09 ORA #IMM 
constant IMORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000010010001"; -- 0x09 ORA #IMM 
constant IMEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010010010000"; -- 0x49 EOR #IMM 
constant IMEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010010010001"; -- 0x49 EOR #IMM 
constant IMCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110010010000"; -- 0xC9 CMP #IMM 
constant IMCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110010010001"; -- 0xC9 CMP #IMM 
constant IMCPX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000000000"; -- 0xE0 CPX #IMM 
constant IMCPX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000000001"; -- 0xE0 CPX #IMM 
constant IMCPY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000000000"; -- 0xC0 CPY #IMM 
constant IMCPY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000000001"; -- 0xC0 CPY #IMM 
constant IMBRK_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010010000"; -- 0x89 BRK #IMM 
constant IMBRK_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010010001"; -- 0x89 BRK #IMM 
constant IMSEP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000100000"; -- 0xE2 SEP #IMM 
constant IMREP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000100000"; -- 0xC2 REP #IMM 
constant IMBIT_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010010000"; -- 0x89 BIT #IMM 
constant IMBIT_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100010010001"; -- 0x89 BIT #IMM 

------------------------------------
--           ZERO PAGE            --
------------------------------------
constant ZPLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001010000"; -- 0xA5 LDA ZP
constant ZPLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001010001"; -- 0xA5 LDA ZP
constant ZPLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001010010"; -- 0xA5 LDA ZP
constant ZPLDX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001100000"; -- 0xA6 LDX ZP
constant ZPLDX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001100001"; -- 0xA6 LDX ZP
constant ZPLDX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001100010"; -- 0xA6 LDX ZP
constant ZPLDY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001000000"; -- 0xA4 LDY ZP
constant ZPLDY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001000001"; -- 0xA4 LDY ZP
constant ZPLDY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001000010"; -- 0xA4 LDY ZP
constant ZPSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001010000"; -- 0x85 STA ZP
constant ZPSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001010001"; -- 0x85 STA ZP
constant ZPSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001010010"; -- 0x85 STA ZP
constant ZPSTX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001100000"; -- 0x86 STX ZP
constant ZPSTX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001100001"; -- 0x86 STX ZP
constant ZPSTX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001100010"; -- 0x86 STX ZP
constant ZPSTY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001000000"; -- 0x84 STY ZP
constant ZPSTY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001000001"; -- 0x84 STY ZP
constant ZPSTY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001000010"; -- 0x84 STY ZP
constant ZPSTZ_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001000000"; -- 0x64 STZ ZP
constant ZPSTZ_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001000001"; -- 0x64 STZ ZP
constant ZPSTZ_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001000010"; -- 0x64 STZ ZP
constant ZPADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001010000"; -- 0x65 ADC ZP
constant ZPADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001010001"; -- 0x65 ADC ZP
constant ZPADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001010010"; -- 0x65 ADC ZP
constant ZPADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001010011"; -- 0x65 ADC ZP
constant ZPSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001010000"; -- 0xE5 SBC ZP
constant ZPSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001010001"; -- 0xE5 SBC ZP
constant ZPSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001010010"; -- 0xE5 SBC ZP
constant ZPSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001010011"; -- 0xE5 SBC ZP
constant ZPCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001010000"; -- 0xC5 CMP ZP
constant ZPCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001010001"; -- 0xC5 CMP ZP
constant ZPCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001010010"; -- 0xC5 CMP ZP
constant ZPCPX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001000000"; -- 0xE4 CPX ZP
constant ZPCPX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001000001"; -- 0xE4 CPX ZP
constant ZPCPX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001000010"; -- 0xE4 CPX ZP
constant ZPCPY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001000000"; -- 0xC4 CPY ZP
constant ZPCPY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001000001"; -- 0xC4 CPY ZP
constant ZPCPY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001000010"; -- 0xC4 CPY ZP
constant ZPAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001010000"; -- 0x25 AND ZP
constant ZPAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001010001"; -- 0x25 AND ZP
constant ZPAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001010010"; -- 0x25 AND ZP
constant ZPORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001010000"; -- 0x05 ORA ZP
constant ZPORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001010001"; -- 0x05 ORA ZP
constant ZPORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001010010"; -- 0x05 ORA ZP
constant ZPEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001010000"; -- 0x45 EOR ZP
constant ZPEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001010001"; -- 0x45 EOR ZP
constant ZPEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001010010"; -- 0x45 EOR ZP
constant ZPBIT_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001000000"; -- 0x24 BIT ZP
constant ZPBIT_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001000001"; -- 0x24 BIT ZP
constant ZPBIT_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001000010"; -- 0x24 BIT ZP
constant ZPASL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001100000"; -- 0x06 ASL ZP 
constant ZPASL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001100001"; -- 0x06 ASL ZP 
constant ZPASL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001100010"; -- 0x06 ASL ZP 
constant ZPASL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001100011"; -- 0x06 ASL ZP 
constant ZPASL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001100100"; -- 0x06 ASL ZP 
constant ZPASL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001100101"; -- 0x06 ASL ZP 
constant ZPLSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001100000"; -- 0x46 LSR ZP 
constant ZPLSR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001100001"; -- 0x46 LSR ZP 
constant ZPLSR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001100010"; -- 0x46 LSR ZP 
constant ZPLSR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001100011"; -- 0x46 LSR ZP 
constant ZPLSR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001100100"; -- 0x46 LSR ZP 
constant ZPLSR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001100101"; -- 0x46 LSR ZP 
constant ZPROL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001100000"; -- 0x26 ROL ZP 
constant ZPROL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001100001"; -- 0x26 ROL ZP 
constant ZPROL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001100010"; -- 0x26 ROL ZP 
constant ZPROL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001100011"; -- 0x26 ROL ZP 
constant ZPROL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001100100"; -- 0x26 ROL ZP 
constant ZPROL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001100101"; -- 0x26 ROL ZP 
constant ZPROR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001100000"; -- 0x66 ROR ZP 
constant ZPROR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001100001"; -- 0x66 ROR ZP 
constant ZPROR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001100010"; -- 0x66 ROR ZP 
constant ZPROR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001100011"; -- 0x66 ROR ZP 
constant ZPROR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001100100"; -- 0x66 ROR ZP 
constant ZPROR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001100101"; -- 0x66 ROR ZP 
constant ZPINC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001100000"; -- 0xE6 INC ZP 
constant ZPINC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001100001"; -- 0xE6 INC ZP 
constant ZPINC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001100010"; -- 0xE6 INC ZP 
constant ZPINC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001100011"; -- 0xE6 INC ZP 
constant ZPINC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001100100"; -- 0xE6 INC ZP 
constant ZPINC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001100101"; -- 0xE6 INC ZP 
constant ZPDEC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001100000"; -- 0xC6 DEC ZP 
constant ZPDEC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001100001"; -- 0xC6 DEC ZP 
constant ZPDEC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001100010"; -- 0xC6 DEC ZP 
constant ZPDEC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001100011"; -- 0xC6 DEC ZP 
constant ZPDEC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001100100"; -- 0xC6 DEC ZP 
constant ZPDEC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001100101"; -- 0xC6 DEC ZP 
constant ZPTSB_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000000"; -- 0x04 TSB ZP 
constant ZPTSB_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000001"; -- 0x04 TSB ZP 
constant ZPTSB_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000010"; -- 0x04 TSB ZP 
constant ZPTSB_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000011"; -- 0x04 TSB ZP 
constant ZPTSB_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000100"; -- 0x04 TSB ZP 
constant ZPTSB_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000101"; -- 0x04 TSB ZP 
constant ZPTSB_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001000110"; -- 0x04 TSB ZP 
constant ZPTRB_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000000"; -- 0x14 TRB ZP 
constant ZPTRB_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000001"; -- 0x14 TRB ZP 
constant ZPTRB_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000010"; -- 0x14 TRB ZP 
constant ZPTRB_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000011"; -- 0x14 TRB ZP 
constant ZPTRB_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000100"; -- 0x14 TRB ZP 
constant ZPTRB_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000101"; -- 0x14 TRB ZP 
constant ZPTRB_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101000110"; -- 0x14 TRB ZP 

------------------------------------
--          ZERO PAGE,X           --
------------------------------------
constant ZXLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101010000"; -- 0xB5 LDA ZP,X
constant ZXLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101010001"; -- 0xB5 LDA ZP,X
constant ZXLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101010010"; -- 0xB5 LDA ZP,X
constant ZXLDY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101000000"; -- 0xB4 LDY ZP,X
constant ZXLDY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101000001"; -- 0xB4 LDY ZP,X
constant ZXLDY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101000010"; -- 0xB4 LDY ZP,X
constant ZXSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101010000"; -- 0x95 STA ZP,X
constant ZXSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101010001"; -- 0x95 STA ZP,X
constant ZXSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101010010"; -- 0x95 STA ZP,X
constant ZXSTY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101000000"; -- 0x94 STY ZP,X
constant ZXSTY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101000001"; -- 0x94 STY ZP,X
constant ZXSTY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101000010"; -- 0x94 STY ZP,X
constant ZXSTZ_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101000000"; -- 0x74 STZ ZP,X
constant ZXSTZ_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101000001"; -- 0x74 STZ ZP,X
constant ZXSTZ_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101000010"; -- 0x74 STZ ZP,X
constant ZXADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101010000"; -- 0x75 ADC ZP,X
constant ZXADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101010001"; -- 0x75 ADC ZP,X
constant ZXADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101010010"; -- 0x75 ADC ZP,X
constant ZXSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101010000"; -- 0xF5 SBC ZP,X
constant ZXSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101010001"; -- 0xF5 SBC ZP,X
constant ZXSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101010010"; -- 0xF5 SBC ZP,X
constant ZXCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101010000"; -- 0xD5 CMP ZP,X
constant ZXCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101010001"; -- 0xD5 CMP ZP,X
constant ZXCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101010010"; -- 0xD5 CMP ZP,X
constant ZXAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101010000"; -- 0x35 AND ZP,X
constant ZXAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101010001"; -- 0x35 AND ZP,X
constant ZXAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101010010"; -- 0x35 AND ZP,X
constant ZXORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101010000"; -- 0x15 ORA ZP,X
constant ZXORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101010001"; -- 0x15 ORA ZP,X
constant ZXORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101010010"; -- 0x15 ORA ZP,X
constant ZXEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101010000"; -- 0x55 EOR ZP,X
constant ZXEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101010001"; -- 0x55 EOR ZP,X
constant ZXEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101010010"; -- 0x55 EOR ZP,X
constant ZXASL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101100000"; -- 0x16 ASL ZP,X
constant ZXASL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101100001"; -- 0x16 ASL ZP,X
constant ZXASL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101100010"; -- 0x16 ASL ZP,X
constant ZXASL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101100011"; -- 0x16 ASL ZP,X
constant ZXASL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101100100"; -- 0x16 ASL ZP,X
constant ZXASL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101100101"; -- 0x16 ASL ZP,X
constant ZXLSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101100000"; -- 0x56 LSR ZP,X
constant ZXLSR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101100001"; -- 0x56 LSR ZP,X
constant ZXLSR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101100010"; -- 0x56 LSR ZP,X
constant ZXLSR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101100011"; -- 0x56 LSR ZP,X
constant ZXLSR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101100100"; -- 0x56 LSR ZP,X
constant ZXLSR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101100101"; -- 0x56 LSR ZP,X
constant ZXROL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101100000"; -- 0x36 ROL ZP,X
constant ZXROL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101100001"; -- 0x36 ROL ZP,X
constant ZXROL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101100010"; -- 0x36 ROL ZP,X
constant ZXROL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101100011"; -- 0x36 ROL ZP,X
constant ZXROL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101100100"; -- 0x36 ROL ZP,X
constant ZXROL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101100101"; -- 0x36 ROL ZP,X
constant ZXROR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101100000"; -- 0x76 ROR ZP,X
constant ZXROR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101100001"; -- 0x76 ROR ZP,X
constant ZXROR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101100010"; -- 0x76 ROR ZP,X
constant ZXROR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101100011"; -- 0x76 ROR ZP,X
constant ZXROR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101100100"; -- 0x76 ROR ZP,X
constant ZXROR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101100101"; -- 0x76 ROR ZP,X
constant ZXDEC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101100000"; -- 0xD6 DEC ZP,X
constant ZXDEC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101100001"; -- 0xD6 DEC ZP,X
constant ZXDEC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101100010"; -- 0xD6 DEC ZP,X
constant ZXDEC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101100011"; -- 0xD6 DEC ZP,X
constant ZXDEC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101100100"; -- 0xD6 DEC ZP,X
constant ZXDEC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101100101"; -- 0xD6 DEC ZP,X
constant ZXINC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101100000"; -- 0xF6 INC ZP,X
constant ZXINC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101100001"; -- 0xF6 INC ZP,X
constant ZXINC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101100010"; -- 0xF6 INC ZP,X
constant ZXINC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101100011"; -- 0xF6 INC ZP,X
constant ZXINC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101100100"; -- 0xF6 INC ZP,X
constant ZXINC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101100101"; -- 0xF6 INC ZP,X
constant ZXBIT_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101000000"; -- 0x34 BIT ZP,X
constant ZXBIT_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101000001"; -- 0x34 BIT ZP,X
constant ZXBIT_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101000010"; -- 0x34 BIT ZP,X

------------------------------------
--          ZERO PAGE,Y           --
------------------------------------
constant ZYLDX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101100000"; -- 0xB6 LDX ZP,Y
constant ZYLDX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101100001"; -- 0xB6 LDX ZP,Y
constant ZYLDX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101100010"; -- 0xB6 LDX ZP,Y
constant ZYLDX_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101100011"; -- 0xB6 LDX ZP,Y

constant ZYSTX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101100000"; -- 0x96 STX ZP,Y
constant ZYSTX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101100001"; -- 0x96 STX ZP,Y
constant ZYSTX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101100010"; -- 0x96 STX ZP,Y

------------------------------------
--           INDIRECT             --
------------------------------------
constant INJMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011000000"; -- 0x6C JMP (IND)
constant INJMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011000001"; -- 0x6C JMP (IND)
constant INJMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011000010"; -- 0x6C JMP (IND)
constant INJMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011000011"; -- 0x6C JMP (IND)
constant INJML_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111000000"; -- 0xDC JML (IND)
constant INJML_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111000001"; -- 0xDC JML (IND)
constant INJML_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111000010"; -- 0xDC JML (IND)
constant INJML_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111000011"; -- 0xDC JML (IND)
constant INJML_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111000100"; -- 0xDC JML (IND)


------------------------------------
--          INDIRECT,Y            --
------------------------------------
constant IYLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100010000"; -- 0xB1 LDA [DIR],Y
constant IYLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100010001"; -- 0xB1 LDA [DIR],Y
constant IYLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100010010"; -- 0xB1 LDA [DIR],Y
constant IYLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100010011"; -- 0xB1 LDA [DIR],Y
constant IYLDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100010100"; -- 0xB1 LDA [DIR],Y
constant IYLDA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100010101"; -- 0xB1 LDA [DIR],Y
constant IYSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100010000"; -- 0x91 STA [DIR],Y
constant IYSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100010001"; -- 0x91 STA [DIR],Y
constant IYSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100010010"; -- 0x91 STA [DIR],Y
constant IYSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100010011"; -- 0x91 STA [DIR],Y
constant IYSTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100010100"; -- 0x91 STA [DIR],Y
constant IYSTA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100010101"; -- 0x91 STA [DIR],Y
constant IYADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100010000"; -- 0x71 ADC [DIR],Y
constant IYADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100010001"; -- 0x71 ADC [DIR],Y
constant IYADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100010010"; -- 0x71 ADC [DIR],Y
constant IYADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100010011"; -- 0x71 ADC [DIR],Y
constant IYADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100010100"; -- 0x71 ADC [DIR],Y
constant IYADC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100010101"; -- 0x71 ADC [DIR],Y
constant IYSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100010000"; -- 0xF1 SBC [DIR],Y
constant IYSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100010001"; -- 0xF1 SBC [DIR],Y
constant IYSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100010010"; -- 0xF1 SBC [DIR],Y
constant IYSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100010011"; -- 0xF1 SBC [DIR],Y
constant IYSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100010100"; -- 0xF1 SBC [DIR],Y
constant IYSBC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100010101"; -- 0xF1 SBC [DIR],Y
constant IYCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100010000"; -- 0xD1 CMP [DIR],Y
constant IYCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100010001"; -- 0xD1 CMP [DIR],Y
constant IYCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100010010"; -- 0xD1 CMP [DIR],Y
constant IYCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100010011"; -- 0xD1 CMP [DIR],Y
constant IYCMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100010100"; -- 0xD1 CMP [DIR],Y
constant IYCMP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100010101"; -- 0xD1 CMP [DIR],Y
constant IYAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100010000"; -- 0x31 AND [DIR],Y
constant IYAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100010001"; -- 0x31 AND [DIR],Y
constant IYAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100010010"; -- 0x31 AND [DIR],Y
constant IYAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100010011"; -- 0x31 AND [DIR],Y
constant IYAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100010100"; -- 0x31 AND [DIR],Y
constant IYAND_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100010101"; -- 0x31 AND [DIR],Y
constant IYORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100010000"; -- 0x11 ORA [DIR],Y
constant IYORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100010001"; -- 0x11 ORA [DIR],Y
constant IYORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100010010"; -- 0x11 ORA [DIR],Y
constant IYORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100010011"; -- 0x11 ORA [DIR],Y
constant IYORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100010100"; -- 0x11 ORA [DIR],Y
constant IYORA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100010101"; -- 0x11 ORA [DIR],Y
constant IYEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100010000"; -- 0x51 EOR [DIR],Y
constant IYEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100010001"; -- 0x51 EOR [DIR],Y
constant IYEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100010010"; -- 0x51 EOR [DIR],Y
constant IYEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100010011"; -- 0x51 EOR [DIR],Y
constant IYEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100010100"; -- 0x51 EOR [DIR],Y
constant IYEOR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100010101"; -- 0x51 EOR [DIR],Y

------------------------------------
--          INDIRECT,X            --
------------------------------------
constant IXLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000010000"; -- 0xA1 LDA (IND_ZP,X)
constant IXLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000010001"; -- 0xA1 LDA (IND_ZP,X)
constant IXLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000010010"; -- 0xA1 LDA (IND_ZP,X)
constant IXLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000010011"; -- 0xA1 LDA (IND_ZP,X)
constant IXLDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000010100"; -- 0xA1 LDA (IND_ZP,X)
constant IXSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000010000"; -- 0x81 STA (IND_ZP,X)
constant IXSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000010001"; -- 0x81 STA (IND_ZP,X)
constant IXSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000010010"; -- 0x81 STA (IND_ZP,X)
constant IXSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000010011"; -- 0x81 STA (IND_ZP,X)
constant IXSTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000010100"; -- 0x81 STA (IND_ZP,X)
constant IXAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000010000"; -- 0x21 AND (IND_ZP,X)
constant IXAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000010001"; -- 0x21 AND (IND_ZP,X)
constant IXAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000010010"; -- 0x21 AND (IND_ZP,X)
constant IXAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000010011"; -- 0x21 AND (IND_ZP,X)
constant IXAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000010100"; -- 0x21 AND (IND_ZP,X)
constant IXORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000010000"; -- 0x01 ORA (IND_ZP,X)
constant IXORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000010001"; -- 0x01 ORA (IND_ZP,X)
constant IXORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000010010"; -- 0x01 ORA (IND_ZP,X)
constant IXORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000010011"; -- 0x01 ORA (IND_ZP,X)
constant IXORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000010100"; -- 0x01 ORA (IND_ZP,X)
constant IXEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000010000"; -- 0x41 EOR (IND_ZP,X)
constant IXEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000010001"; -- 0x41 EOR (IND_ZP,X)
constant IXEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000010010"; -- 0x41 EOR (IND_ZP,X)
constant IXEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000010011"; -- 0x41 EOR (IND_ZP,X)
constant IXEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000010100"; -- 0x41 EOR (IND_ZP,X)
constant IXCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000010000"; -- 0xC1 CMP (IND_ZP,X)
constant IXCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000010001"; -- 0xC1 CMP (IND_ZP,X)
constant IXCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000010010"; -- 0xC1 CMP (IND_ZP,X)
constant IXCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000010011"; -- 0xC1 CMP (IND_ZP,X)
constant IXCMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000010100"; -- 0xC1 CMP (IND_ZP,X)
constant IXADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000010000"; -- 0x61 ADC (IND_ZP,X)
constant IXADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000010001"; -- 0x61 ADC (IND_ZP,X)
constant IXADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000010010"; -- 0x61 ADC (IND_ZP,X)
constant IXADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000010011"; -- 0x61 ADC (IND_ZP,X)
constant IXADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000010100"; -- 0x61 ADC (IND_ZP,X)
constant IXSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000010000"; -- 0xE1 SBC (IND_ZP,X)
constant IXSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000010001"; -- 0xE1 SBC (IND_ZP,X)
constant IXSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000010010"; -- 0xE1 SBC (IND_ZP,X)
constant IXSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000010011"; -- 0xE1 SBC (IND_ZP,X)
constant IXSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000010100"; -- 0xE1 SBC (IND_ZP,X)
constant IXJMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111000000"; -- 0x7C JMP (IND,X)
constant IXJMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111000001"; -- 0x7C JMP (IND,X)
constant IXJMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111000010"; -- 0x7C JMP (IND,X)
constant IXJMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111000011"; -- 0x7C JMP (IND,X)
constant IXJMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111000100"; -- 0x7C JMP (IND,X)
constant IXJSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111000000"; -- 0xFC JSR (IND,X)
constant IXJSR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111000001"; -- 0xFC JSR (IND,X)
constant IXJSR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111000010"; -- 0xFC JSR (IND,X)
constant IXJSR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111000011"; -- 0xFC JSR (IND,X)
constant IXJSR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111000100"; -- 0xFC JSR (IND,X)
constant IXJSR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111000101"; -- 0xFC JSR (IND,X)

------------------------------------
--            ABSOLUTE            --
------------------------------------
constant ABLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011010000"; -- 0xAD LDA ABS
constant ABLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011010001"; -- 0xAD LDA ABS
constant ABLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011010010"; -- 0xAD LDA ABS
constant ABLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011010011"; -- 0xAD LDA ABS
constant ABLDX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011100000"; -- 0xAE LDX ABS
constant ABLDX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011100001"; -- 0xAE LDX ABS
constant ABLDX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011100010"; -- 0xAE LDX ABS
constant ABLDX_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011100011"; -- 0xAE LDX ABS
constant ABLDY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011000000"; -- 0xAC LDY ABS
constant ABLDY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011000001"; -- 0xAC LDY ABS
constant ABLDY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011000010"; -- 0xAC LDY ABS
constant ABLDY_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011000011"; -- 0xAC LDY ABS
constant ABSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011010000"; -- 0x8D STA ABS
constant ABSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011010001"; -- 0x8D STA ABS
constant ABSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011010010"; -- 0x8D STA ABS
constant ABSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011010011"; -- 0x8D STA ABS
constant ABSTX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011100000"; -- 0x8E STX ABS
constant ABSTX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011100001"; -- 0x8E STX ABS
constant ABSTX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011100010"; -- 0x8E STX ABS
constant ABSTX_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011100011"; -- 0x8E STX ABS
constant ABSTY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011000000"; -- 0x8C STY ABS
constant ABSTY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011000001"; -- 0x8C STY ABS
constant ABSTY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011000010"; -- 0x8C STY ABS
constant ABSTY_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011000011"; -- 0x8C STY ABS
constant ABSTZ_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111000000"; -- 0x9C STZ ABS
constant ABSTZ_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111000001"; -- 0x9C STZ ABS
constant ABSTZ_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111000010"; -- 0x9C STZ ABS
constant ABSTZ_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111000011"; -- 0x9C STZ ABS
constant ABADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011010000"; -- 0x6D ADC ABS
constant ABADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011010001"; -- 0x6D ADC ABS
constant ABADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011010010"; -- 0x6D ADC ABS
constant ABADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011010011"; -- 0x6D ADC ABS
constant ABADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011010100"; -- 0x6D ADC ABS
constant ABSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011010000"; -- 0xED SBC ABS
constant ABSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011010001"; -- 0xED SBC ABS
constant ABSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011010010"; -- 0xED SBC ABS
constant ABSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011010011"; -- 0xED SBC ABS
constant ABSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011010100"; -- 0xED SBC ABS
constant ABORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011010000"; -- 0x0D ORA ABS
constant ABORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011010001"; -- 0x0D ORA ABS
constant ABORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011010010"; -- 0x0D ORA ABS
constant ABORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011010011"; -- 0x0D ORA ABS
constant ABAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011010000"; -- 0x2D AND ABS
constant ABAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011010001"; -- 0x2D AND ABS
constant ABAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011010010"; -- 0x2D AND ABS
constant ABAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011010011"; -- 0x2D AND ABS
constant ABEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011010000"; -- 0x4D EOR ABS
constant ABEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011010001"; -- 0x4D EOR ABS
constant ABEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011010010"; -- 0x4D EOR ABS
constant ABEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011010011"; -- 0x4D EOR ABS
constant ABCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011010000"; -- 0xCD CMP ABS
constant ABCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011010001"; -- 0xCD CMP ABS
constant ABCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011010010"; -- 0xCD CMP ABS
constant ABCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011010011"; -- 0xCD CMP ABS
constant ABCPX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011000000"; -- 0xEC CPX ABS
constant ABCPX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011000001"; -- 0xEC CPX ABS
constant ABCPX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011000010"; -- 0xEC CPX ABS
constant ABCPX_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011000011"; -- 0xEC CPX ABS
constant ABCPY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011000000"; -- 0xCC CPY ABS
constant ABCPY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011000001"; -- 0xCC CPY ABS
constant ABCPY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011000010"; -- 0xCC CPY ABS
constant ABCPY_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011000011"; -- 0xCC CPY ABS
constant ABJMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011000000"; -- 0x4C JMP ABS
constant ABJMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011000001"; -- 0x4C JMP ABS
constant ABJSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000000000"; -- 0x20 JSR ABS
constant ABJSR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000000001"; -- 0x20 JSR ABS
constant ABJSR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000000010"; -- 0x20 JSR ABS
constant ABJSR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000000011"; -- 0x20 JSR ABS
constant ABBIT_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011000000"; -- 0x2C BIT ABS
constant ABBIT_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011000001"; -- 0x2C BIT ABS
constant ABBIT_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011000010"; -- 0x2C BIT ABS
constant ABBIT_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011000011"; -- 0x2C BIT ABS
constant ABASL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100000"; -- 0x0E ASL ABS
constant ABASL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100001"; -- 0x0E ASL ABS
constant ABASL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100010"; -- 0x0E ASL ABS
constant ABASL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100011"; -- 0x0E ASL ABS
constant ABASL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100100"; -- 0x0E ASL ABS
constant ABASL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100101"; -- 0x0E ASL ABS
constant ABASL_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011100110"; -- 0x0E ASL ABS
constant ABLSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100000"; -- 0x4E LSR ABS
constant ABLSR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100001"; -- 0x4E LSR ABS
constant ABLSR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100010"; -- 0x4E LSR ABS
constant ABLSR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100011"; -- 0x4E LSR ABS
constant ABLSR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100100"; -- 0x4E LSR ABS
constant ABLSR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100101"; -- 0x4E LSR ABS
constant ABLSR_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011100110"; -- 0x4E LSR ABS
constant ABROL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100000"; -- 0x2E ROL ABS
constant ABROL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100001"; -- 0x2E ROL ABS
constant ABROL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100010"; -- 0x2E ROL ABS
constant ABROL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100011"; -- 0x2E ROL ABS
constant ABROL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100100"; -- 0x2E ROL ABS
constant ABROL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100101"; -- 0x2E ROL ABS
constant ABROL_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011100110"; -- 0x2E ROL ABS
constant ABROR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100000"; -- 0x6E ROR ABS
constant ABROR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100001"; -- 0x6E ROR ABS
constant ABROR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100010"; -- 0x6E ROR ABS
constant ABROR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100011"; -- 0x6E ROR ABS
constant ABROR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100100"; -- 0x6E ROR ABS
constant ABROR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100101"; -- 0x6E ROR ABS
constant ABROR_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011100110"; -- 0x6E ROR ABS
constant ABINC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100000"; -- 0xEE INC ABS
constant ABINC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100001"; -- 0xEE INC ABS
constant ABINC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100010"; -- 0xEE INC ABS
constant ABINC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100011"; -- 0xEE INC ABS
constant ABINC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100100"; -- 0xEE INC ABS
constant ABINC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100101"; -- 0xEE INC ABS
constant ABINC_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011100110"; -- 0xEE INC ABS
constant ABDEC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100000"; -- 0xCE DEC ABS
constant ABDEC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100001"; -- 0xCE DEC ABS
constant ABDEC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100010"; -- 0xCE DEC ABS
constant ABDEC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100011"; -- 0xCE DEC ABS
constant ABDEC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100100"; -- 0xCE DEC ABS
constant ABDEC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100101"; -- 0xCE DEC ABS
constant ABDEC_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011100110"; -- 0xCE DEC ABS
constant ABTSB_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000000"; -- 0x0C TSB ABS
constant ABTSB_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000001"; -- 0x0C TSB ABS
constant ABTSB_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000010"; -- 0x0C TSB ABS
constant ABTSB_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000011"; -- 0x0C TSB ABS
constant ABTSB_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000100"; -- 0x0C TSB ABS
constant ABTSB_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000101"; -- 0x0C TSB ABS
constant ABTSB_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000110"; -- 0x0C TSB ABS
constant ABTSB_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011000111"; -- 0x0C TSB ABS
constant ABTRB_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000000"; -- 0x1C TRB ABS
constant ABTRB_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000001"; -- 0x1C TRB ABS
constant ABTRB_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000010"; -- 0x1C TRB ABS
constant ABTRB_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000011"; -- 0x1C TRB ABS
constant ABTRB_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000100"; -- 0x1C TRB ABS
constant ABTRB_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000101"; -- 0x1C TRB ABS
constant ABTRB_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000110"; -- 0x1C TRB ABS
constant ABTRB_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111000111"; -- 0x1C TRB ABS

------------------------------------
--           ABSOLUTE,X           --
------------------------------------
constant AXLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111010000"; -- 0xBD LDA ABS,X
constant AXLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111010001"; -- 0xBD LDA ABS,X
constant AXLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111010010"; -- 0xBD LDA ABS,X
constant AXLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111010011"; -- 0xBD LDA ABS,X
constant AXLDY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111000000"; -- 0xBC LDY ABS,X
constant AXLDY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111000001"; -- 0xBC LDY ABS,X
constant AXLDY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111000010"; -- 0xBC LDY ABS,X
constant AXLDY_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111000011"; -- 0xBC LDY ABS,X
constant AXSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111010000"; -- 0x9D STA ABS,X
constant AXSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111010001"; -- 0x9D STA ABS,X
constant AXSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111010010"; -- 0x9D STA ABS,X
constant AXSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111010011"; -- 0x9D STA ABS,X
constant AXSTZ_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111100000"; -- 0x9E STZ ABS,X
constant AXSTZ_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111100001"; -- 0x9E STZ ABS,X
constant AXSTZ_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111100010"; -- 0x9E STZ ABS,X
constant AXSTZ_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111100011"; -- 0x9E STZ ABS,X
constant AXADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111010000"; -- 0x7D ADC ABS,X
constant AXADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111010001"; -- 0x7D ADC ABS,X
constant AXADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111010010"; -- 0x7D ADC ABS,X
constant AXADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111010011"; -- 0x7D ADC ABS,X
constant AXSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111010000"; -- 0xFD SBC ABS,X
constant AXSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111010001"; -- 0xFD SBC ABS,X
constant AXSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111010010"; -- 0xFD SBC ABS,X
constant AXSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111010011"; -- 0xFD SBC ABS,X
constant AXCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111010000"; -- 0xDD CMP ABS,X
constant AXCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111010001"; -- 0xDD CMP ABS,X
constant AXCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111010010"; -- 0xDD CMP ABS,X
constant AXCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111010011"; -- 0xDD CMP ABS,X
constant AXINC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100000"; -- 0xFE INC ABS,X
constant AXINC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100001"; -- 0xFE INC ABS,X
constant AXINC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100010"; -- 0xFE INC ABS,X
constant AXINC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100011"; -- 0xFE INC ABS,X
constant AXINC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100100"; -- 0xFE INC ABS,X
constant AXINC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100101"; -- 0xFE INC ABS,X
constant AXINC_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111100110"; -- 0xFE INC ABS,X
constant AXDEC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100000"; -- 0xDE DEC ABS,X
constant AXDEC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100001"; -- 0xDE DEC ABS,X
constant AXDEC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100010"; -- 0xDE DEC ABS,X
constant AXDEC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100011"; -- 0xDE DEC ABS,X
constant AXDEC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100100"; -- 0xDE DEC ABS,X
constant AXDEC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100101"; -- 0xDE DEC ABS,X
constant AXDEC_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111100110"; -- 0xDE DEC ABS,X
constant AXASL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100000"; -- 0x1E ASL ABS,X
constant AXASL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100001"; -- 0x1E ASL ABS,X
constant AXASL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100010"; -- 0x1E ASL ABS,X
constant AXASL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100011"; -- 0x1E ASL ABS,X
constant AXASL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100100"; -- 0x1E ASL ABS,X
constant AXASL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100101"; -- 0x1E ASL ABS,X
constant AXASL_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111100110"; -- 0x1E ASL ABS,X
constant AXLSR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100000"; -- 0x5E LSR ABS,X
constant AXLSR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100001"; -- 0x5E LSR ABS,X
constant AXLSR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100010"; -- 0x5E LSR ABS,X
constant AXLSR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100011"; -- 0x5E LSR ABS,X
constant AXLSR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100100"; -- 0x5E LSR ABS,X
constant AXLSR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100101"; -- 0x5E LSR ABS,X
constant AXLSR_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111100110"; -- 0x5E LSR ABS,X
constant AXROL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100000"; -- 0x3E ROL ABS,X
constant AXROL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100001"; -- 0x3E ROL ABS,X
constant AXROL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100010"; -- 0x3E ROL ABS,X
constant AXROL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100011"; -- 0x3E ROL ABS,X
constant AXROL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100100"; -- 0x3E ROL ABS,X
constant AXROL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100101"; -- 0x3E ROL ABS,X
constant AXROL_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111100110"; -- 0x3E ROL ABS,X
constant AXROR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100000"; -- 0x7E ROR ABS,X
constant AXROR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100001"; -- 0x7E ROR ABS,X
constant AXROR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100010"; -- 0x7E ROR ABS,X
constant AXROR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100011"; -- 0x7E ROR ABS,X
constant AXROR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100100"; -- 0x7E ROR ABS,X
constant AXROR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100101"; -- 0x7E ROR ABS,X
constant AXROR_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111100110"; -- 0x7E ROR ABS,X
constant AXAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111010000"; -- 0x3D AND ABS,X
constant AXAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111010001"; -- 0x3D AND ABS,X
constant AXAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111010010"; -- 0x3D AND ABS,X
constant AXAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111010011"; -- 0x3D AND ABS,X
constant AXORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111010000"; -- 0x1D ORA ABS,X
constant AXORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111010001"; -- 0x1D ORA ABS,X
constant AXORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111010010"; -- 0x1D ORA ABS,X
constant AXORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111010011"; -- 0x1D ORA ABS,X
constant AXEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111010000"; -- 0x5D EOR ABS,X
constant AXEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111010001"; -- 0x5D EOR ABS,X
constant AXEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111010010"; -- 0x5D EOR ABS,X
constant AXEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111010011"; -- 0x5D EOR ABS,X
constant AXBIT_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111000000"; -- 0x3C BIT ABS,X
constant AXBIT_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111000001"; -- 0x3C BIT ABS,X
constant AXBIT_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111000010"; -- 0x3C BIT ABS,X
constant AXBIT_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111000011"; -- 0x3C BIT ABS,X

------------------------------------
--           ABSOLUTE,Y           --
------------------------------------
constant AYLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110010000"; -- 0xB9 LDA ABS,Y
constant AYLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110010001"; -- 0xB9 LDA ABS,Y
constant AYLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110010010"; -- 0xB9 LDA ABS,Y
constant AYLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101110010011"; -- 0xB9 LDA ABS,Y
constant AYLDX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111100000"; -- 0xBE LDX ABS,Y
constant AYLDX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111100001"; -- 0xBE LDX ABS,Y
constant AYLDX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111100010"; -- 0xBE LDX ABS,Y
constant AYLDX_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111100011"; -- 0xBE LDX ABS,Y
constant AYSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110010000"; -- 0x99 STA ABS,Y
constant AYSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110010001"; -- 0x99 STA ABS,Y
constant AYSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110010010"; -- 0x99 STA ABS,Y
constant AYSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100110010011"; -- 0x99 STA ABS,Y
constant AYADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110010000"; -- 0x79 ADC ABS,Y
constant AYADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110010001"; -- 0x79 ADC ABS,Y
constant AYADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110010010"; -- 0x79 ADC ABS,Y
constant AYADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110010011"; -- 0x79 ADC ABS,Y
constant AYADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011110010100"; -- 0x79 ADC ABS,Y
constant AYSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110010000"; -- 0xF9 SBC ABS,Y
constant AYSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110010001"; -- 0xF9 SBC ABS,Y
constant AYSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110010010"; -- 0xF9 SBC ABS,Y
constant AYSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110010011"; -- 0xF9 SBC ABS,Y
constant AYSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111110010100"; -- 0xF9 SBC ABS,Y
constant AYCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110010000"; -- 0xD9 CMP ABS,Y
constant AYCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110010001"; -- 0xD9 CMP ABS,Y
constant AYCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110010010"; -- 0xD9 CMP ABS,Y
constant AYCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110110010011"; -- 0xD9 CMP ABS,Y
constant AYORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110010000"; -- 0x19 ORA ABS,Y
constant AYORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110010001"; -- 0x19 ORA ABS,Y
constant AYORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110010010"; -- 0x19 ORA ABS,Y
constant AYORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000110010011"; -- 0x19 ORA ABS,Y
constant AYAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110010000"; -- 0x39 AND ABS,Y
constant AYAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110010001"; -- 0x39 AND ABS,Y
constant AYAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110010010"; -- 0x39 AND ABS,Y
constant AYAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001110010011"; -- 0x39 AND ABS,Y
constant AYEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110010000"; -- 0x59 EOR ABS,Y
constant AYEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110010001"; -- 0x59 EOR ABS,Y
constant AYEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110010010"; -- 0x59 EOR ABS,Y
constant AYEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010110010011"; -- 0x59 EOR ABS,Y

------------------------------------------------
--           ABSOLUTE LONG (JUMP...)          --
------------------------------------------------
constant ABJML_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111000000"; -- 0x5C JML ABS
constant ABJML_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111000001"; -- 0x5C JML ABS
constant ABJML_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111000010"; -- 0x5C JML ABS
constant ABJSL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000100000"; -- 0x22 JSL ABS
constant ABJSL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000100001"; -- 0x22 JSL ABS
constant ABJSL_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000100010"; -- 0x22 JSL ABS
constant ABJSL_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000100011"; -- 0x22 JSL ABS
constant ABJSL_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000100100"; -- 0x22 JSL ABS
constant ABJSL_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000100101"; -- 0x22 JSL ABS

------------------------------------
--           RELATIVE             --
------------------------------------
constant   BRA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000000000"; -- 0x80 BRA       
constant   BCC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100000000"; -- 0x90 BCC       
constant   BCS_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100000000"; -- 0xB0 BCS       
constant   BEQ_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100000000"; -- 0xF0 BEQ       
constant   BNE_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100000000"; -- 0xD0 BNE       
constant   BPL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100000000"; -- 0x10 BPL       
constant   BMI_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100000000"; -- 0x30 BMI       
constant   BVC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100000000"; -- 0x50 BVC       
constant   BVS_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100000000"; -- 0x70 BVS       

---------------------------------------
--           RELATIVE LONG           --
---------------------------------------
constant   BRL_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000100000"; -- 0x82 BRL       
constant   BRL_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000100001"; -- 0x82 BRL       

-------------------------------
--           STACK           --
-------------------------------
constant   PEA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101000000"; -- 0xF4 PEA
constant   PEA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101000001"; -- 0xF4 PEA
constant   PEA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101000010"; -- 0xF4 PEA
constant   PEA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101000011"; -- 0xF4 PEA
constant   PEI_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101000000"; -- 0xD4 PEI
constant   PEI_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101000001"; -- 0xD4 PEI
constant   PEI_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101000010"; -- 0xD4 PEI
constant   PEI_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101000011"; -- 0xD4 PEI
constant   PEI_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101000100"; -- 0xD4 PEI
constant   PER_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000100000"; -- 0x62 PER
constant   PER_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000100001"; -- 0x62 PER
constant   PER_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000100010"; -- 0x62 PER
constant   PER_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000100011"; -- 0x62 PER
constant   PER_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000100100"; -- 0x62 PER

----------------------------------
--          DIRECT,Y            --
----------------------------------
constant DYLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110000"; -- 0xB7 LDA [DIR],Y
constant DYLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110001"; -- 0xB7 LDA [DIR],Y
constant DYLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110010"; -- 0xB7 LDA [IND],Y
constant DYLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110011"; -- 0xB7 LDA [DIR],Y
constant DYLDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110100"; -- 0xB7 LDA [DIR],Y
constant DYLDA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110101"; -- 0xB7 LDA [DIR],Y
constant DYLDA_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101101110110"; -- 0xB7 LDA [DIR],Y
constant DYSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110000"; -- 0x97 STA [DIR],Y
constant DYSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110001"; -- 0x97 STA [DIR],Y
constant DYSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110010"; -- 0x97 STA [DIR],Y
constant DYSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110011"; -- 0x97 STA [DIR],Y
constant DYSTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110100"; -- 0x97 STA [DIR],Y
constant DYSTA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110101"; -- 0x97 STA [DIR],Y
constant DYSTA_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100101110110"; -- 0x97 STA [DIR],Y
constant DYADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110000"; -- 0x77 ADC [DIR],Y
constant DYADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110001"; -- 0x77 ADC [DIR],Y
constant DYADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110010"; -- 0x77 ADC [DIR],Y
constant DYADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110011"; -- 0x77 ADC [DIR],Y
constant DYADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110100"; -- 0x77 ADC [DIR],Y
constant DYADC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110101"; -- 0x77 ADC [DIR],Y
constant DYADC_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011101110110"; -- 0x77 ADC [DIR],Y
constant DYSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110000"; -- 0xF7 SBC [DIR],Y
constant DYSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110001"; -- 0xF7 SBC [DIR],Y
constant DYSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110010"; -- 0xF7 SBC [DIR],Y
constant DYSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110011"; -- 0xF7 SBC [DIR],Y
constant DYSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110100"; -- 0xF7 SBC [DIR],Y
constant DYSBC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110101"; -- 0xF7 SBC [DIR],Y
constant DYSBC_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111101110110"; -- 0xF7 SBC [DIR],Y
constant DYCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110000"; -- 0xD7 CMP [DIR],Y
constant DYCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110001"; -- 0xD7 CMP [DIR],Y
constant DYCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110010"; -- 0xD7 CMP [DIR],Y
constant DYCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110011"; -- 0xD7 CMP [DIR],Y
constant DYCMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110100"; -- 0xD7 CMP [DIR],Y
constant DYCMP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110101"; -- 0xD7 CMP [DIR],Y
constant DYCMP_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110101110110"; -- 0xD7 CMP [DIR],Y
constant DYAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110000"; -- 0x37 AND [DIR],Y
constant DYAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110001"; -- 0x37 AND [DIR],Y
constant DYAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110010"; -- 0x37 AND [DIR],Y
constant DYAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110011"; -- 0x37 AND [DIR],Y
constant DYAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110100"; -- 0x37 AND [DIR],Y
constant DYAND_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110101"; -- 0x37 AND [DIR],Y
constant DYAND_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001101110110"; -- 0x37 AND [DIR],Y
constant DYORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110000"; -- 0x17 ORA [DIR],Y
constant DYORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110001"; -- 0x17 ORA [DIR],Y
constant DYORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110010"; -- 0x17 ORA [DIR],Y
constant DYORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110011"; -- 0x17 ORA [DIR],Y
constant DYORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110100"; -- 0x17 ORA [DIR],Y
constant DYORA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110101"; -- 0x17 ORA [DIR],Y
constant DYORA_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000101110110"; -- 0x17 ORA [DIR],Y
constant DYEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110000"; -- 0x57 EOR [DIR],Y
constant DYEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110001"; -- 0x57 EOR [DIR],Y
constant DYEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110010"; -- 0x57 EOR [DIR],Y
constant DYEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110011"; -- 0x57 EOR [DIR],Y
constant DYEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110100"; -- 0x57 EOR [DIR],Y
constant DYEOR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110101"; -- 0x57 EOR [DIR],Y
constant DYEOR_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101110110"; -- 0x57 EOR [DIR],Y

--------------------------------
--          DIRECT            --
--------------------------------
constant DILDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001110000"; -- 0xA7 LDA [DIR]
constant DILDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001110001"; -- 0xA7 LDA [DIR]
constant DILDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001110010"; -- 0xA7 LDA [IND]
constant DILDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001110011"; -- 0xA7 LDA [DIR]
constant DILDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001110100"; -- 0xA7 LDA [DIR]
constant DILDA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101001110101"; -- 0xA7 LDA [DIR]
constant DISTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001110000"; -- 0x87 STA [DIR]
constant DISTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001110001"; -- 0x87 STA [DIR]
constant DISTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001110010"; -- 0x87 STA [DIR]
constant DISTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001110011"; -- 0x87 STA [DIR]
constant DISTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001110100"; -- 0x87 STA [DIR]
constant DISTA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100001110101"; -- 0x87 STA [DIR]
constant DIADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001110000"; -- 0x67 ADC [DIR]
constant DIADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001110001"; -- 0x67 ADC [DIR]
constant DIADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001110010"; -- 0x67 ADC [DIR]
constant DIADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001110011"; -- 0x67 ADC [DIR]
constant DIADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001110100"; -- 0x67 ADC [DIR]
constant DIADC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011001110101"; -- 0x67 ADC [DIR]
constant DISBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001110000"; -- 0xE7 SBC [DIR]
constant DISBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001110001"; -- 0xE7 SBC [DIR]
constant DISBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001110010"; -- 0xE7 SBC [DIR]
constant DISBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001110011"; -- 0xE7 SBC [DIR]
constant DISBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001110100"; -- 0xE7 SBC [DIR]
constant DISBC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111001110101"; -- 0xE7 SBC [DIR]
constant DICMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001110000"; -- 0xC7 CMP [DIR]
constant DICMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001110001"; -- 0xC7 CMP [DIR]
constant DICMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001110010"; -- 0xC7 CMP [DIR]
constant DICMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001110011"; -- 0xC7 CMP [DIR]
constant DICMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001110100"; -- 0xC7 CMP [DIR]
constant DICMP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110001110101"; -- 0xC7 CMP [DIR]
constant DIAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001110000"; -- 0x27 AND [DIR]
constant DIAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001110001"; -- 0x27 AND [DIR]
constant DIAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001110010"; -- 0x27 AND [DIR]
constant DIAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001110011"; -- 0x27 AND [DIR]
constant DIAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001110100"; -- 0x27 AND [DIR]
constant DIAND_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001001110101"; -- 0x27 AND [DIR]
constant DIORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001110000"; -- 0x07 ORA [DIR]
constant DIORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001110001"; -- 0x07 ORA [DIR]
constant DIORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001110010"; -- 0x07 ORA [DIR]
constant DIORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001110011"; -- 0x07 ORA [DIR]
constant DIORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001110100"; -- 0x07 ORA [DIR]
constant DIORA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000001110101"; -- 0x07 ORA [DIR]
constant DIEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001110000"; -- 0x47 EOR [DIR]
constant DIEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001110001"; -- 0x47 EOR [DIR]
constant DIEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001110010"; -- 0x47 EOR [DIR]
constant DIEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001110011"; -- 0x47 EOR [DIR]
constant DIEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001110100"; -- 0x47 EOR [DIR]
constant DIEOR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001110101"; -- 0x47 EOR [DIR]

----------------------------------------
--            ABSOLUTE LONG           --
----------------------------------------
constant ALLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011110000"; -- 0xAF LDA ABS_LONG
constant ALLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011110001"; -- 0xAF LDA ABS_LONG
constant ALLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011110010"; -- 0xAF LDA ABS_LONG
constant ALLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011110011"; -- 0xAF LDA ABS_LONG
constant ALLDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101011110100"; -- 0xAF LDA ABS_LONG
constant ALSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011110000"; -- 0x8F STA ABS_LONG
constant ALSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011110001"; -- 0x8F STA ABS_LONG
constant ALSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011110010"; -- 0x8F STA ABS_LONG
constant ALSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011110011"; -- 0x8F STA ABS_LONG
constant ALSTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100011110100"; -- 0x8F STA ABS_LONG
constant ALADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011110000"; -- 0x6F ADC ABS_LONG
constant ALADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011110001"; -- 0x6F ADC ABS_LONG
constant ALADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011110010"; -- 0x6F ADC ABS_LONG
constant ALADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011110011"; -- 0x6F ADC ABS_LONG
constant ALADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011110100"; -- 0x6F ADC ABS_LONG
constant ALADC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011011110101"; -- 0x6F ADC ABS_LONG
constant ALSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011110000"; -- 0xEF SBC ABS_LONG
constant ALSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011110001"; -- 0xEF SBC ABS_LONG
constant ALSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011110010"; -- 0xEF SBC ABS_LONG
constant ALSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011110011"; -- 0xEF SBC ABS_LONG
constant ALSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011110100"; -- 0xEF SBC ABS_LONG
constant ALSBC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111011110101"; -- 0xEF SBC ABS_LONG
constant ALORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011110000"; -- 0x0F ORA ABS_LONG
constant ALORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011110001"; -- 0x0F ORA ABS_LONG
constant ALORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011110010"; -- 0x0F ORA ABS_LONG
constant ALORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011110011"; -- 0x0F ORA ABS_LONG
constant ALORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000011110100"; -- 0x0F ORA ABS_LONG
constant ALAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011110000"; -- 0x2F AND ABS_LONG
constant ALAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011110001"; -- 0x2F AND ABS_LONG
constant ALAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011110010"; -- 0x2F AND ABS_LONG
constant ALAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011110011"; -- 0x2F AND ABS_LONG
constant ALAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001011110100"; -- 0x2F AND ABS_LONG
constant ALEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011110000"; -- 0x4F EOR ABS_LONG
constant ALEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011110001"; -- 0x4F EOR ABS_LONG
constant ALEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011110010"; -- 0x4F EOR ABS_LONG
constant ALEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011110011"; -- 0x4F EOR ABS_LONG
constant ALEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010011110100"; -- 0x4F EOR ABS_LONG
constant ALCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011110000"; -- 0xCF CMP ABS_LONG
constant ALCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011110001"; -- 0xCF CMP ABS_LONG
constant ALCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011110010"; -- 0xCF CMP ABS_LONG
constant ALCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011110011"; -- 0xCF CMP ABS_LONG
constant ALCMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110011110100"; -- 0xCF CMP ABS_LONG

-----------------------------------------
--           ABSOLUTE LONG,X           --
-----------------------------------------
constant AILDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111110000"; -- 0xBF LDA ABS_LONG,X
constant AILDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111110001"; -- 0xBF LDA ABS_LONG,X
constant AILDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111110010"; -- 0xBF LDA ABS_LONG,X
constant AILDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111110011"; -- 0xBF LDA ABS_LONG,X
constant AILDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111110100"; -- 0xBF LDA ABS_LONG,X
constant AILDA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101111110101"; -- 0xBF LDA ABS_LONG,X
constant AISTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111110000"; -- 0x9F STA ABS_LONG,X
constant AISTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111110001"; -- 0x9F STA ABS_LONG,X
constant AISTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111110010"; -- 0x9F STA ABS_LONG,X
constant AISTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111110011"; -- 0x9F STA ABS_LONG,X
constant AISTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111110100"; -- 0x9F STA ABS_LONG,X
constant AISTA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100111110101"; -- 0x9F STA ABS_LONG,X
constant AIADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111110000"; -- 0x7F ADC ABS_LONG,X
constant AIADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111110001"; -- 0x7F ADC ABS_LONG,X
constant AIADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111110010"; -- 0x7F ADC ABS_LONG,X
constant AIADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111110011"; -- 0x7F ADC ABS_LONG,X
constant AIADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111110100"; -- 0x7F ADC ABS_LONG,X
constant AIADC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011111110101"; -- 0x7F ADC ABS_LONG,X
constant AISBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111110000"; -- 0xFF SBC ABS_LONG,X
constant AISBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111110001"; -- 0xFF SBC ABS_LONG,X
constant AISBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111110010"; -- 0xFF SBC ABS_LONG,X
constant AISBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111110011"; -- 0xFF SBC ABS_LONG,X
constant AISBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111110100"; -- 0xFF SBC ABS_LONG,X
constant AISBC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111111110101"; -- 0xFF SBC ABS_LONG,X
constant AICMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111110000"; -- 0xDF CMP ABS_LONG,X
constant AICMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111110001"; -- 0xDF CMP ABS_LONG,X
constant AICMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111110010"; -- 0xDF CMP ABS_LONG,X
constant AICMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111110011"; -- 0xDF CMP ABS_LONG,X
constant AICMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111110100"; -- 0xDF CMP ABS_LONG,X
constant AICMP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110111110101"; -- 0xDF CMP ABS_LONG,X
constant AIAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111110000"; -- 0x3F AND ABS_LONG,X
constant AIAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111110001"; -- 0x3F AND ABS_LONG,X
constant AIAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111110010"; -- 0x3F AND ABS_LONG,X
constant AIAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111110011"; -- 0x3F AND ABS_LONG,X
constant AIAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111110100"; -- 0x3F AND ABS_LONG,X
constant AIAND_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001111110101"; -- 0x3F AND ABS_LONG,X
constant AIORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111110000"; -- 0x1F ORA ABS_LONG,X
constant AIORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111110001"; -- 0x1F ORA ABS_LONG,X
constant AIORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111110010"; -- 0x1F ORA ABS_LONG,X
constant AIORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111110011"; -- 0x1F ORA ABS_LONG,X
constant AIORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111110100"; -- 0x1F ORA ABS_LONG,X
constant AIORA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000111110101"; -- 0x1F ORA ABS_LONG,X
constant AIEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111110000"; -- 0x5F EOR ABS_LONG,X
constant AIEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111110001"; -- 0x5F EOR ABS_LONG,X
constant AIEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111110010"; -- 0x5F EOR ABS_LONG,X
constant AIEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111110011"; -- 0x5F EOR ABS_LONG,X
constant AIEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111110100"; -- 0x5F EOR ABS_LONG,X
constant AIEOR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010111110101"; -- 0x5F EOR ABS_LONG,X

-----------------------------------------
--            STACK RELATIVE           --
-----------------------------------------
constant SRLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000110000"; -- 0xA3 LDA $XX,S
constant SRLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000110001"; -- 0xA3 LDA $XX,S
constant SRLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101000110010"; -- 0xA3 LDA $XX,S
constant SRSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000110000"; -- 0x83 STA $XX,S
constant SRSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000110001"; -- 0x83 STA $XX,S
constant SRSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100000110010"; -- 0x83 STA $XX,S
constant SRADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000110000"; -- 0x63 ADC $XX,S
constant SRADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000110001"; -- 0x63 ADC $XX,S
constant SRADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011000110010"; -- 0x63 ADC $XX,S
constant SRSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000110000"; -- 0xE3 SBC $XX,S
constant SRSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000110001"; -- 0xE3 SBC $XX,S
constant SRSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111000110010"; -- 0xE3 SBC $XX,S
constant SRCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000110000"; -- 0xC3 CMP $XX,S
constant SRCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000110001"; -- 0xC3 CMP $XX,S
constant SRCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110000110010"; -- 0xC3 CMP $XX,S
constant SRAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000110000"; -- 0x23 AND $XX,S
constant SRAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000110001"; -- 0x23 AND $XX,S
constant SRAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001000110010"; -- 0x23 AND $XX,S
constant SRORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000110000"; -- 0x03 ORA $XX,S
constant SRORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000110001"; -- 0x03 ORA $XX,S
constant SRORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000000110010"; -- 0x03 ORA $XX,S
constant SREOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000110000"; -- 0x43 EOR $XX,S
constant SREOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000110001"; -- 0x43 EOR $XX,S
constant SREOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010000110010"; -- 0x43 EOR $XX,S

--------------------------------------------------
--            STACK RELATIVE INDEXED Y          --
--------------------------------------------------
constant SYLDA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100110000"; -- 0xB3 LDA ($XX,S),Y
constant SYLDA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100110001"; -- 0xB3 LDA ($XX,S),Y
constant SYLDA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100110010"; -- 0xB3 LDA ($XX,S),Y
constant SYLDA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100110011"; -- 0xB3 LDA ($XX,S),Y
constant SYLDA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100110100"; -- 0xB3 LDA ($XX,S),Y
constant SYLDA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0101100110101"; -- 0xB3 LDA ($XX,S),Y
constant SYSTA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100110000"; -- 0x93 STA ($XX,S),Y
constant SYSTA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100110001"; -- 0x93 STA ($XX,S),Y
constant SYSTA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100110010"; -- 0x93 STA ($XX,S),Y
constant SYSTA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100110011"; -- 0x93 STA ($XX,S),Y
constant SYSTA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100110100"; -- 0x93 STA ($XX,S),Y
constant SYSTA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0100100110101"; -- 0x93 STA ($XX,S),Y
constant SYADC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100110000"; -- 0x73 ADC ($XX,S),Y
constant SYADC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100110001"; -- 0x73 ADC ($XX,S),Y
constant SYADC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100110010"; -- 0x73 ADC ($XX,S),Y
constant SYADC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100110011"; -- 0x73 ADC ($XX,S),Y
constant SYADC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100110100"; -- 0x73 ADC ($XX,S),Y
constant SYADC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0011100110101"; -- 0x73 ADC ($XX,S),Y
constant SYSBC_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100110000"; -- 0xF3 SBC ($XX,S),Y
constant SYSBC_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100110001"; -- 0xF3 SBC ($XX,S),Y
constant SYSBC_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100110010"; -- 0xF3 SBC ($XX,S),Y
constant SYSBC_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100110011"; -- 0xF3 SBC ($XX,S),Y
constant SYSBC_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100110100"; -- 0xF3 SBC ($XX,S),Y
constant SYSBC_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0111100110101"; -- 0xF3 SBC ($XX,S),Y
constant SYCMP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100110000"; -- 0xD3 CMP ($XX,S),Y
constant SYCMP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100110001"; -- 0xD3 CMP ($XX,S),Y
constant SYCMP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100110010"; -- 0xD3 CMP ($XX,S),Y
constant SYCMP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100110011"; -- 0xD3 CMP ($XX,S),Y
constant SYCMP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100110100"; -- 0xD3 CMP ($XX,S),Y
constant SYCMP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0110100110101"; -- 0xD3 CMP ($XX,S),Y
constant SYAND_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100110000"; -- 0x33 AND ($XX,S),Y
constant SYAND_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100110001"; -- 0x33 AND ($XX,S),Y
constant SYAND_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100110010"; -- 0x33 AND ($XX,S),Y
constant SYAND_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100110011"; -- 0x33 AND ($XX,S),Y
constant SYAND_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100110100"; -- 0x33 AND ($XX,S),Y
constant SYAND_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0001100110101"; -- 0x33 AND ($XX,S),Y
constant SYORA_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100110000"; -- 0x13 ORA ($XX,S),Y
constant SYORA_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100110001"; -- 0x13 ORA ($XX,S),Y
constant SYORA_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100110010"; -- 0x13 ORA ($XX,S),Y
constant SYORA_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100110011"; -- 0x13 ORA ($XX,S),Y
constant SYORA_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100110100"; -- 0x13 ORA ($XX,S),Y
constant SYORA_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0000100110101"; -- 0x13 ORA ($XX,S),Y
constant SYEOR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100110000"; -- 0x53 EOR ($XX,S),Y
constant SYEOR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100110001"; -- 0x53 EOR ($XX,S),Y
constant SYEOR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100110010"; -- 0x53 EOR ($XX,S),Y
constant SYEOR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100110011"; -- 0x53 EOR ($XX,S),Y
constant SYEOR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100110100"; -- 0x53 EOR ($XX,S),Y
constant SYEOR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010100110101"; -- 0x53 EOR ($XX,S),Y

------------------------------------
--           MOVE BLOCK           --
------------------------------------
constant MBMVN_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000000"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000001"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000010"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000011"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000100"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000101"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000110"; -- 0x54 MVN $xx,$xx
constant MBMVN_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010101000111"; -- 0x54 MVN $xx,$xx

constant MBMVP_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000000"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000001"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000010"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000011"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000100"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000101"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000110"; -- 0x44 MVP $xx,$xx
constant MBMVP_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "0010001000111"; -- 0x44 MVP $xx,$xx

-------------------------------------------------
--           NEW OPCODES (WDM OPCODE)          --
-------------------------------------------------
-- IMPLIED
constant   PHR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100010110000"; -- 0x8B PHR AXY->S (two byte instruction)
constant   PHR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100010110001"; -- 0x8B PHR AXY->S (two byte instruction)
constant   PHR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100010110010"; -- 0x8B PHR AXY->S (two byte instruction)
constant   PHR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100010110011"; -- 0x8B PHR AXY->S (two byte instruction)
constant   PHR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100010110100"; -- 0x8B PHR AXY->S (two byte instruction)
constant   PHR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100010110101"; -- 0x8B PHR AXY->S (two byte instruction)

constant   PLR_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110000"; -- 0xAB PLR S->YXA (two byte instruction)
constant   PLR_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110001"; -- 0xAB PLR S->YXA (two byte instruction)
constant   PLR_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110010"; -- 0xAB PLR S->YXA (two byte instruction)
constant   PLR_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110011"; -- 0xAB PLR S->YXA (two byte instruction)
constant   PLR_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110100"; -- 0xAB PLR S->YXA (two byte instruction)
constant   PLR_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110101"; -- 0xAB PLR S->YXA (two byte instruction)
constant   PLR_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1101010110110"; -- 0xAB PLR S->YXA (two byte instruction)

constant   SAV_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000000"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000001"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000010"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000011"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000100"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000101"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000110"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100000111"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP8: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100001000"; -- 0x90 SAV AXYBDP->S (two byte instruction)
constant   SAV_OP9: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100001001"; -- 0x90 SAV AXYBDP->S (two byte instruction)

constant   RST_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010000"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010001"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010010"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010011"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP4: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010100"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP5: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010101"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP6: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010110"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP7: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100010111"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP8: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100011000"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant   RST_OP9: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100011001"; -- 0x91 RST S->PDBYXA (two byte instruction)
constant  RST_OP10: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100100011010"; -- 0x91 RST S->PDBYXA (two byte instruction)

-- MULTIPLY UNSIGNED 16X16->32 BIT
constant   MPU_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011100000"; -- 0x8E MPU multiply A*X (two byte instruction)
constant   MPU_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011100001"; -- 0x8E MPU multiply A*X (two byte instruction)
constant   MPU_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011100010"; -- 0x8E MPU multiply A*X (two byte instruction)
constant   MPU_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011100011"; -- 0x8E MPU multiply A*X (two byte instruction)

-- MULTIPLY SIGNED 16X16->32 BIT
constant   MPS_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011110000"; -- 0x8F MPS multiply A*X (two byte instruction)
constant   MPS_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011110001"; -- 0x8F MPS multiply A*X (two byte instruction)
constant   MPS_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011110010"; -- 0x8F MPS multiply A*X (two byte instruction)
constant   MPS_OP3: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1100011110011"; -- 0x8F MPS multiply A*X (two byte instruction)

-- REGISTERS EXCHANGE
constant   XYX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1111010110000"; -- 0xEB EXCHANGE X <-> Y (two byte instruction)
constant   XYX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1111010110001"; -- 0xEB EXCHANGE X <-> Y (two byte instruction)
constant   XYX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1111010110010"; -- 0xEB EXCHANGE X <-> Y (two byte instruction)
constant   XAX_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1000010110000"; -- 0x0B EXCHANGE A <-> X (two byte instruction)
constant   XAX_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1000010110001"; -- 0x0B EXCHANGE A <-> X (two byte instruction)
constant   XAX_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1000010110010"; -- 0x0B EXCHANGE A <-> X (two byte instruction)
constant   XAY_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1001010110000"; -- 0x2B EXCHANGE A <-> Y (two byte instruction)
constant   XAY_OP1: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1001010110001"; -- 0x2B EXCHANGE A <-> Y (two byte instruction)
constant   XAY_OP2: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1001010110010"; -- 0x2B EXCHANGE A <-> Y (two byte instruction)

-- MISC
constant   EXT_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1111011000000"; -- 0xEC EXTEND SIGN OF A TO B (two byte instruction)
constant   NEG_OP0: STD_LOGIC_VECTOR(MC_ADDR_LENGTH downto 0) :=  "1111011010000"; -- 0xED NEGATE A         (two byte instruction)

 
-- ALU microcode
constant NOP_A: STD_LOGIC_VECTOR(4 downto 0) := "00000";    -- no operation
constant SUM_A: STD_LOGIC_VECTOR(4 downto 0) := "00001";    -- sum with carry
constant SUB_A: STD_LOGIC_VECTOR(4 downto 0) := "00010";    -- subtract with borrow
constant AND_A: STD_LOGIC_VECTOR(4 downto 0) := "00011";    -- and
constant  OR_A: STD_LOGIC_VECTOR(4 downto 0) := "00100";    -- or
constant XOR_A: STD_LOGIC_VECTOR(4 downto 0) := "00101";    -- xor
constant INC_A: STD_LOGIC_VECTOR(4 downto 0) := "00110";    -- increment by 1
constant DEC_A: STD_LOGIC_VECTOR(4 downto 0) := "00111";    -- decrement by 1
constant SHL_A: STD_LOGIC_VECTOR(4 downto 0) := "01000";    -- shift left
constant SHR_A: STD_LOGIC_VECTOR(4 downto 0) := "01001";    -- shift right
constant ROL_A: STD_LOGIC_VECTOR(4 downto 0) := "01010";    -- rotation left
constant ROR_A: STD_LOGIC_VECTOR(4 downto 0) := "01011";    -- rotation right
constant SWC_A: STD_LOGIC_VECTOR(4 downto 0) := "01100";    -- sum without carry (used for indexing and branches)
constant SWC_N: STD_LOGIC_VECTOR(4 downto 0) := "01100";    -- subtract without borrow (used only by branches with negative offset)
constant BIT_A: STD_LOGIC_VECTOR(4 downto 0) := "01101";    -- bit test (used by BIT opcode)
constant DAA_A: STD_LOGIC_VECTOR(4 downto 0) := "01110";    -- decimal adjustement for BCD sum
constant DAS_A: STD_LOGIC_VECTOR(4 downto 0) := "01111";    -- decimal adjustement for BCD subtract
constant CMP_A: STD_LOGIC_VECTOR(4 downto 0) := "10000";    -- compare
constant TSB_A: STD_LOGIC_VECTOR(4 downto 0) := "10001";    -- test and set bit
constant TRB_A: STD_LOGIC_VECTOR(4 downto 0) := "10010";    -- test and reset bit
constant EXT_A: STD_LOGIC_VECTOR(4 downto 0) := "10011";    -- extend sign
constant NEG_A: STD_LOGIC_VECTOR(4 downto 0) := "10100";    -- negate

-- PCR microcode
constant NOP_PC: STD_LOGIC_VECTOR(3 downto 0) := "0000"; -- PC no operation
constant LSB_PC: STD_LOGIC_VECTOR(3 downto 0) := "0001"; -- PC load lsb
constant MSB_PC: STD_LOGIC_VECTOR(3 downto 0) := "0010"; -- PC load msb
constant INC_PC: STD_LOGIC_VECTOR(3 downto 0) := "0011"; -- PC increment by 1
constant LOD_PC: STD_LOGIC_VECTOR(3 downto 0) := "0100"; -- PC load lsb\msb  (used by JMP\JSR instructions)
constant LML_PC: STD_LOGIC_VECTOR(3 downto 0) := "0101"; -- PC load lsb\msb from oper register (used for JML\JSL instructions)
constant IN2_PC: STD_LOGIC_VECTOR(3 downto 0) := "0110"; -- PC = PC +2 (BRK opcode)
constant DE3_PC: STD_LOGIC_VECTOR(3 downto 0) := "0111"; -- PC = PC -3 (MVN/MVP opcodes)
constant BRA_PC: STD_LOGIC_VECTOR(3 downto 0) := "1000"; -- PC branch
constant BRL_PC: STD_LOGIC_VECTOR(3 downto 0) := "1001"; -- PC branch long 

-- MPR (memory data pointer) microcode
constant NOP_M: STD_LOGIC_VECTOR(4 downto 0) := "00000"; -- no operation
constant LSB_M: STD_LOGIC_VECTOR(4 downto 0) := "00001"; -- load lsb
constant MSB_M: STD_LOGIC_VECTOR(4 downto 0) := "00010"; -- load msb
constant INC_M: STD_LOGIC_VECTOR(4 downto 0) := "00011"; -- increment 
constant DEC_M: STD_LOGIC_VECTOR(4 downto 0) := "00100"; -- decrement
constant VEC_M: STD_LOGIC_VECTOR(4 downto 0) := "00101"; -- load vector
constant ZPL_M: STD_LOGIC_VECTOR(4 downto 0) := "00110"; -- load ZEROPAGE
constant ALL_M: STD_LOGIC_VECTOR(4 downto 0) := "00111"; -- load all 16 bit register
constant ICC_M: STD_LOGIC_VECTOR(4 downto 0) := "01000"; -- increment MSB with carry
constant DOX_M: STD_LOGIC_VECTOR(4 downto 0) := "01001"; -- add D + offset + X
constant DOY_M: STD_LOGIC_VECTOR(4 downto 0) := "01010"; -- add D + offset + Y
constant AOS_M: STD_LOGIC_VECTOR(4 downto 0) := "01011"; -- add S + offset
constant ABX_M: STD_LOGIC_VECTOR(4 downto 0) := "01100"; -- add opr+X
constant ABY_M: STD_LOGIC_VECTOR(4 downto 0) := "01101"; -- add opr+Y
constant ADX_M: STD_LOGIC_VECTOR(4 downto 0) := "01110"; -- add X
constant ADY_M: STD_LOGIC_VECTOR(4 downto 0) := "01111"; -- add Y
constant MHB_M: STD_LOGIC_VECTOR(4 downto 0) := "10000"; -- load high byte 
constant AOY_M: STD_LOGIC_VECTOR(4 downto 0) := "10001"; -- add opr+Y and concatenates SBR

-- address multiplexer microcode
constant ADPC: STD_LOGIC_VECTOR(2 downto 0) := "000";  -- select PC
constant ADMP: STD_LOGIC_VECTOR(2 downto 0) := "001";  -- select MP
constant ADSP: STD_LOGIC_VECTOR(2 downto 0) := "010";  -- select SP
constant ADDI: STD_LOGIC_VECTOR(2 downto 0) := "011";  -- select Direct
constant ADXR: STD_LOGIC_VECTOR(2 downto 0) := "100";  -- select X register
constant ADYR: STD_LOGIC_VECTOR(2 downto 0) := "101";  -- select Y register
constant ADNP: STD_LOGIC_VECTOR(2 downto 0) := "000";  -- no operation (PC)

-- PR microcode
constant NOP_P: STD_LOGIC_VECTOR(4 downto 0) := "00000"; -- PR no operation
constant PLD_P: STD_LOGIC_VECTOR(4 downto 0) := "00001"; -- PR load
constant FLD_P: STD_LOGIC_VECTOR(4 downto 0) := "00010"; -- NV load
constant FLC_P: STD_LOGIC_VECTOR(4 downto 0) := "00011"; -- NZC load
constant FLV_P: STD_LOGIC_VECTOR(4 downto 0) := "00100"; -- NVZC load
constant SEC_P: STD_LOGIC_VECTOR(4 downto 0) := "00101"; -- 1 => C 
constant CLC_P: STD_LOGIC_VECTOR(4 downto 0) := "00110"; -- 0 => C 
constant SEI_P: STD_LOGIC_VECTOR(4 downto 0) := "00111"; -- 1 => I 
constant CLI_P: STD_LOGIC_VECTOR(4 downto 0) := "01000"; -- 0 => I 
constant SED_P: STD_LOGIC_VECTOR(4 downto 0) := "01001"; -- 1 => D 
constant CLD_P: STD_LOGIC_VECTOR(4 downto 0) := "01010"; -- 0 => D 
constant CLV_P: STD_LOGIC_VECTOR(4 downto 0) := "01011"; -- 0 => V 
constant AUC_P: STD_LOGIC_VECTOR(4 downto 0) := "01100"; -- auc => ACR 
constant HAC_P: STD_LOGIC_VECTOR(4 downto 0) := "01101"; -- hold ACR 
constant SID_P: STD_LOGIC_VECTOR(4 downto 0) := "01110"; -- 1 => I/D 
constant LDZ_P: STD_LOGIC_VECTOR(4 downto 0) := "01111"; -- Z load
constant XCE_P: STD_LOGIC_VECTOR(4 downto 0) := "10000"; -- E => C; C => E
constant SEP_P: STD_LOGIC_VECTOR(4 downto 0) := "10001"; -- P = P OR din
constant REP_P: STD_LOGIC_VECTOR(4 downto 0) := "10010"; -- P = P AND not din
constant WDM_P: STD_LOGIC_VECTOR(4 downto 0) := "10011"; -- 1 => op_exp;
constant WDC_P: STD_LOGIC_VECTOR(4 downto 0) := "10100"; -- 0 => op_exp;
constant FLW_P: STD_LOGIC_VECTOR(4 downto 0) := "10101"; -- NZ load, 0 -> op_exp
constant MUF_P: STD_LOGIC_VECTOR(4 downto 0) := "10110"; -- Z load from unsigned multplier
constant MSF_P: STD_LOGIC_VECTOR(4 downto 0) := "10111"; -- NZ load from unsigned multplier

-- register operation microcode REGOP (decreg)
constant NOP_R: STD_LOGIC_VECTOR(5 downto 0) := "000000";  -- no operation
constant ALL_R: STD_LOGIC_VECTOR(5 downto 0) := "000001";  -- register A load lsb
constant ALM_R: STD_LOGIC_VECTOR(5 downto 0) := "000010";  -- register A load msb
constant A16_R: STD_LOGIC_VECTOR(5 downto 0) := "000011";  -- register A load msb & lsb
constant XLL_R: STD_LOGIC_VECTOR(5 downto 0) := "000100";  -- register X load lsb
constant XLM_R: STD_LOGIC_VECTOR(5 downto 0) := "000101";  -- register X load msb 
constant X16_R: STD_LOGIC_VECTOR(5 downto 0) := "000110";  -- register X load msb & lsb 
constant YLL_R: STD_LOGIC_VECTOR(5 downto 0) := "000111";  -- register Y load lsb
constant YLM_R: STD_LOGIC_VECTOR(5 downto 0) := "001000";  -- register Y load msb
constant Y16_R: STD_LOGIC_VECTOR(5 downto 0) := "001001";  -- register Y load msb & lsb
constant DLL_R: STD_LOGIC_VECTOR(5 downto 0) := "001010";  -- register D load lsb
constant DLM_R: STD_LOGIC_VECTOR(5 downto 0) := "001011";  -- register D load msb
constant D16_R: STD_LOGIC_VECTOR(5 downto 0) := "001100";  -- register D load msb & lsb
constant OLD_R: STD_LOGIC_VECTOR(5 downto 0) := "001101";  -- register O load lsb
constant OMD_R: STD_LOGIC_VECTOR(5 downto 0) := "001110";  -- register O load msb
constant SLD_R: STD_LOGIC_VECTOR(5 downto 0) := "001111";  -- register S load lsb
constant SLM_R: STD_LOGIC_VECTOR(5 downto 0) := "010000";  -- register S load msb
constant S16_R: STD_LOGIC_VECTOR(5 downto 0) := "010001";  -- register S load msb & lsb
constant SUP_R: STD_LOGIC_VECTOR(5 downto 0) := "010010";  -- register S increment by 1
constant SDW_R: STD_LOGIC_VECTOR(5 downto 0) := "010011";  -- register S decrement by 1
constant SAU_R: STD_LOGIC_VECTOR(5 downto 0) := "010100";  -- register A (lsb) load/register S increment by 1
constant SXU_R: STD_LOGIC_VECTOR(5 downto 0) := "010101";  -- register X (lsb) load/register S increment by 1
constant SXM_R: STD_LOGIC_VECTOR(5 downto 0) := "010110";  -- register X (msb) load/register S increment by 1
constant SYU_R: STD_LOGIC_VECTOR(5 downto 0) := "010111";  -- register Y (lsb) load/register S increment by 1
constant SYM_R: STD_LOGIC_VECTOR(5 downto 0) := "011000";  -- register Y (msb) load/register S increment by 1
constant KLD_R: STD_LOGIC_VECTOR(5 downto 0) := "011001";  -- register K (PBR) load
constant BLD_R: STD_LOGIC_VECTOR(5 downto 0) := "011010";  -- register B (DBR) load
constant KCL_R: STD_LOGIC_VECTOR(5 downto 0) := "011011";  -- register K (PBR) clear and register S decrement by 1
constant BCL_R: STD_LOGIC_VECTOR(5 downto 0) := "011100";  -- register B (DBR) clear
constant SKC_R: STD_LOGIC_VECTOR(5 downto 0) := "011101";  -- register B (DBR) clear and register S decrement by 1
constant DEA_R: STD_LOGIC_VECTOR(5 downto 0) := "011110";  -- register A decrement (MVN/MVP)
constant O16_R: STD_LOGIC_VECTOR(5 downto 0) := "011111";  -- register O load msb & lsb
constant OSU_R: STD_LOGIC_VECTOR(5 downto 0) := "100000";  -- register O load lsb/register S increment by 1
constant MVN_R: STD_LOGIC_VECTOR(5 downto 0) := "100001";  -- register XY increment by 1, A decremented by 1
constant MVP_R: STD_LOGIC_VECTOR(5 downto 0) := "100010";  -- register XY decrement by 1, A decremented by 1
constant MUL_R: STD_LOGIC_VECTOR(5 downto 0) := "100011";  -- register A/B load multiplication lsb result, register X load multiplication msb result
constant MUI_R: STD_LOGIC_VECTOR(5 downto 0) := "100100";  -- multiplication init
constant MUS_R: STD_LOGIC_VECTOR(5 downto 0) := "100101";  -- multiplication (unsigned) start
constant MSS_R: STD_LOGIC_VECTOR(5 downto 0) := "100110";  -- multiplication (signed) start
constant WAI_R: STD_LOGIC_VECTOR(5 downto 0) := "100111";  -- WAI set flipflop
constant STP_R: STD_LOGIC_VECTOR(5 downto 0) := "101000";  -- STP set flipflop
constant BLS_R: STD_LOGIC_VECTOR(5 downto 0) := "101001";  -- register B (DBR) load/register S incremented by 1
constant DLS_R: STD_LOGIC_VECTOR(5 downto 0) := "101010";  -- register D load msb & lsb/register S incremented by 1

-- register multiplexer microcode RSEL (ALU operand #1)
constant EXT_O: STD_LOGIC_VECTOR(4 downto 0) := "00000";  -- external data bus
constant ARD_O: STD_LOGIC_VECTOR(4 downto 0) := "00001";  -- register A msb & lsb select
constant ARM_O: STD_LOGIC_VECTOR(4 downto 0) := "00010";  -- register A msb select (also returns A swapped)
constant XRD_O: STD_LOGIC_VECTOR(4 downto 0) := "00011";  -- register X msb & lsb select
constant XRM_O: STD_LOGIC_VECTOR(4 downto 0) := "00100";  -- register X msb select
constant YRD_O: STD_LOGIC_VECTOR(4 downto 0) := "00101";  -- register Y msb & lsb select
constant YRM_O: STD_LOGIC_VECTOR(4 downto 0) := "00110";  -- register Y msb select
constant SRD_O: STD_LOGIC_VECTOR(4 downto 0) := "00111";  -- register S lsb select
constant PRD_O: STD_LOGIC_VECTOR(4 downto 0) := "01000";  -- register P select
constant PLR_O: STD_LOGIC_VECTOR(4 downto 0) := "01001";  -- register PCL select
constant PHR_O: STD_LOGIC_VECTOR(4 downto 0) := "01010";  -- register PCH select
constant ORD_O: STD_LOGIC_VECTOR(4 downto 0) := "01011";  -- register O msb & lsb select 
constant Z00_O: STD_LOGIC_VECTOR(4 downto 0) := "01100";  -- select (all zero output)
constant DRD_O: STD_LOGIC_VECTOR(4 downto 0) := "01101";  -- register D msb & lsb select
constant DRM_O: STD_LOGIC_VECTOR(4 downto 0) := "01110";  -- register D msb select
constant KRD_O: STD_LOGIC_VECTOR(4 downto 0) := "01111";  -- register K PBR
constant BRD_O: STD_LOGIC_VECTOR(4 downto 0) := "10000";  -- register B PBR
constant EXM_O: STD_LOGIC_VECTOR(4 downto 0) := "10001";  -- external data bus on MSB, O on lsb
constant OMD_O: STD_LOGIC_VECTOR(4 downto 0) := "10010";  -- register O msb select 
constant PCR_O: STD_LOGIC_VECTOR(4 downto 0) := "10011";  -- register PC (16 bit) select

-- data multiplexer microcode DMUX (ALU operand #2)
constant NOP_D: STD_LOGIC_VECTOR(2 downto 0) := "000";
constant ORD_D: STD_LOGIC_VECTOR(2 downto 0) := "001";
constant EXT_D: STD_LOGIC_VECTOR(2 downto 0) := "010";
constant EXM_D: STD_LOGIC_VECTOR(2 downto 0) := "011";
constant BCD_D: STD_LOGIC_VECTOR(2 downto 0) := "100";

-- read/write control
constant   RDE: STD_LOGIC_VECTOR(1 downto 0) := "11";    -- data bus read
constant   WRE: STD_LOGIC_VECTOR(1 downto 0) := "10";    -- data bus write (combinatorial mode)
constant   WRL: STD_LOGIC_VECTOR(1 downto 0) := "01";    -- data bus write (registered mode)

begin
  process(em,m,x,a)
  begin            
	 -----------------------------------
	 --          NATIVE MODE          --
	 -----------------------------------
    if em = '0' then  
	  -- The PLA is arranged like an ROM, there are an address input "a" and an data output "q". The address of PLA is 13 bit wide 
	  -- and composed in this way:
	  --
	  --  W  ----  CPU OPCODE   ---- --- MPC --
	  --  |  |                     | |        |  
	  --  |  |                     | |        |  
	  --  W  X--X--X--X--X--X--X--X--Y--Y--Y--Y 
	  -- 12-11-10-09-08-07-06-05-04-03-02-01-00
	  --
	  -- the bit (12) W is the two byte instruction bit
	  -- the bits (11-4) (X field) is formed by CPU instruction opcode 
	  -- the bits (3-0) (Y field) is formed by the three bit wide microinstruction program counter (MPC)  
	  -- The MPC field is cleared at each opcode fetch by FSM and since it's three bit wide there are
	  -- an maximum of eight microinstructions available per opcode 
	  --
	  -- The bits 10-3 of PLA address serves to select the microcode group of a related CPU opcode 
	  -- and they are stable for all instruction execution time, instead the remaining three bit 2-0 (MPC field) of PLA address 
	  -- increment at each clock in order to address the next microcode instructions.   
	  -- microcode assembly:
	  -- Due the particulary pipeline structure of this CPU, all microinstructions have an extra cycle hidden on fetch 
	  -- of the next opcode instruction and normally this extra cycle is coded as "NOP" (see the last line  "when  others =>...").
	  -- However there are some instructions where this extra cycle is used for some functions like decimal adjustments etc of
	  -- ADC and SBC instructions (see DAA and DAS).
	  --
	  -- Microcode fields:
	  --     
	  --                          DMUX: ALU operand #2 multiplexer
	  --                          |       AI: effective address is indexed (X or Y)
	  --                          |       |   VP: vector pull
	  --                          |       |   |   ML: memory lock            
	  --                          |       |   |   |   VPA: valid program address 
	  --                          |       |   |   |   |   VDA: valid data address 
	  --                          |       |   |   |   |   |   EI: end of microcode sequence (the hidden extra cycle it's always executed after this microinstruction) 
	  --                          |       |   |   |   |   |   |   W: read/write control
	  --                          |       |   |   |   |   |   |   |    CLI: clear interrupt request
	  --                          |       |   |   |   |   |   |   |    |    PD: PC/MP address output multiplexer select
	  --                          |       |   |   |   |   |   |   |    |    |      PCR: register PC (program counter)
	  --                          |       |   |   |   |   |   |   |    |    |      |        MPR: register MP (memory pointer)
	  --                          |       |   |   |   |   |   |   |    |    |      |        |       P_OP: register P set/reset bit
	  --                          |       |   |   |   |   |   |   |    |    |      |        |       |       ALUOP: ALU operation
	  --                          |       |   |   |   |   |   |   |    |    |      |        |       |       |       REGOP: registers load/increment/decrement etc.
	  --                          |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       RSEL: registers output multiplexer select
	  --                          |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
	  --                          |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
		 case a is              -- DMUX    AI  VP  ML VPA VDA  EI  W    CLI  PD     PCR      MPR     P_OP    ALUOP   REGOP   RSEL
			------------------------------------
			--            IMPLIED             --
			------------------------------------
			-- BRK
			when    BRK_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & IN2_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- if no interrupt request then PC=PC+2 
			when    BRK_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & KRD_O; -- PBR->S; SP-1 
			when    BRK_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1 
			when    BRK_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1 
			when    BRK_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & VEC_M & SID_P & NOP_A & KCL_R & PRD_O; -- P->S; VEC->MP; CLI; SEI; CLD
			when    BRK_OP5 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'0'& RDE &'1'& ADMP & LSB_PC & INC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCL; MP+1; 1->B; VP
			when    BRK_OP6 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'1'& RDE &'1'& ADMP & MSB_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCH; EI; VP 

			-- COP
			when    COP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & IN2_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- if no interrupt request then PC=PC+2 
			when    COP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & KRD_O; -- PBR->S; SP-1 
			when    COP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1 
			when    COP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1 
			when    COP_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & VEC_M & SID_P & NOP_A & KCL_R & PRD_O; -- P->S; VEC->MP; CLI; SEI; CLD
			when    COP_OP5 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'0'& RDE &'1'& ADMP & LSB_PC & INC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCL; MP+1; 1->B; VP
			when    COP_OP6 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'1'& RDE &'1'& ADMP & MSB_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCH; EI; VP 
			
			-- NOP
		   when    NOP_OP0 => q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- EI
			
			-- CLC
			when    CLC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLC_P & NOP_A & NOP_R & EXT_O; -- 0->C; EI

			-- SEC
			when    SEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & SEC_P & NOP_A & NOP_R & EXT_O; -- 1->C; EI

			-- CLI
			when    CLI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLI_P & NOP_A & NOP_R & EXT_O; -- 0->I; EI

			-- SEI
			when    SEI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & SEI_P & NOP_A & NOP_R & EXT_O; -- 1->I; EI

			-- CLV
			when    CLV_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLV_P & NOP_A & NOP_R & EXT_O; -- 0->V; EI
			
			-- CLD
			when    CLD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLD_P & NOP_A & NOP_R & EXT_O; -- 0->D; EI

			-- SED
			when    SED_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & SED_P & NOP_A & NOP_R & EXT_O; -- 1->D; EI

			-- TAX
			when    TAX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & ARD_O; -- A->X; EI

			-- TXA
			when    TXA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & XRD_O; -- X->A; EI

			-- TAY
			when    TAY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & ARD_O; -- A->Y; EI

			-- TYA
			when    TYA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & YRD_O; -- Y->A; EI

			-- TXY
			when    TXY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & XRD_O; -- X->Y; EI

			-- TYX
			when    TYX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & YRD_O; -- Y->X; EI

			-- TCD
			when    TCD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & D16_R & ARD_O; -- C->D; EI

			-- TDC
			when    TDC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & DRD_O; -- D->C; EI

			-- TXS
			when    TXS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & S16_R & XRD_O; -- X->S; EI

			-- TSX
			when    TSX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & SRD_O; -- S->X; EI

			-- INC A
			when    INC_OP0 => 
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & ALL_R & ARD_O; -- A+1; EI
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & A16_R & ARD_O; -- A+1; EI
                 end if;					  

			-- DEC A
			when    DEC_OP0 => 
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & ALL_R & ARD_O; -- A-1; EI
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & A16_R & ARD_O; -- A-1; EI
                 end if;					  
			
			-- INX
			when    INX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & X16_R & XRD_O; -- X+1; EI

			-- DEX
			when    DEX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & X16_R & XRD_O; -- X-1; EI
			
			-- INY
			when    INY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & Y16_R & YRD_O; -- Y+1; EI

			-- DEY
			when    DEY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & Y16_R & YRD_O; -- Y-1; EI

			-- PHP
			when    PHP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PRD_O; -- P->S; SP-1; EI 

			-- PHD
			when    PHD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & DRM_O; -- D (msb) ->S; SP-1;
			when    PHD_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & DRD_O; -- D (lsb) ->S; SP-1; EI 
			
			-- PHA
			when    PHA_OP0 =>
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A (lsb) ->S; SP-1; EI 
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARM_O; -- A (msb) ->S; SP-1;
               end if;					
			when    PHA_OP1 =>
					if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A (lsb) ->S; SP-1; EI 
               end if;
					
			-- PHX
			when    PHX_OP0 =>
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X (lsb) ->S; SP-1; EI 
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRM_O; -- X (msb) ->S; SP-1;
               end if;					
			when    PHX_OP1 =>
					if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X (lsb) ->S; SP-1; EI 
               end if;

			-- PHY
			when    PHY_OP0 =>
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRD_O; -- Y (lsb) ->S; SP-1; EI 
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRM_O; -- Y (msb) ->S; SP-1;
               end if;					
			when    PHY_OP1 =>
					if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRD_O; -- Y (lsb) ->S; SP-1; EI 
               end if;

			-- PHR (in native mode PHR pushes ALWAYS 16 bit registers)
			when    PHR_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARM_O; -- A(msb)->S; SP-1;     (two byte instruction) 
			when    PHR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A(lsb)->S; SP-1;     (two byte instruction) 
			when    PHR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRM_O; -- X(msb)->S; SP-1;     (two byte instruction)
			when    PHR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X(lsb)->S; SP-1;     (two byte instruction)
			when    PHR_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRM_O; -- Y(msb)->S; SP-1;     (two byte instruction)
			when    PHR_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & SDW_R & YRD_O; -- Y(lsb)->S; SP-1; EI  (two byte instruction)

			-- SAV (in native mode STO pushes ALWAYS AXY 16 bit registers)
			when    SAV_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARM_O; -- A(msb)->S; SP-1;     (two byte instruction) 
			when    SAV_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A(lsb)->S; SP-1;     (two byte instruction) 
			when    SAV_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRM_O; -- X(msb)->S; SP-1;     (two byte instruction)
			when    SAV_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X(lsb)->S; SP-1;     (two byte instruction)
			when    SAV_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRM_O; -- Y(msb)->S; SP-1;     (two byte instruction)
			when    SAV_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRD_O; -- Y(lsb)->S; SP-1;     (two byte instruction)
			when    SAV_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PRD_O; -- P->S; SP-1;          (two byte instruction)
			when    SAV_OP7 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & BRD_O; -- B->S; SP-1;          (two byte instruction)
			when    SAV_OP8 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & DRM_O; -- D (msb) ->S; SP-1;   (two byte instruction)
			when    SAV_OP9 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & SDW_R & DRD_O; -- D (lsb) ->S; SP-1;   (two byte instruction)

			-- RST (in native mode RST pulls ALWAYS AXY 16 bit registers)
			when    RST_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP;     SP+1 (two byte instruction)
			when    RST_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- S->O (lsb); SP+1
			when    RST_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & DLS_R & EXM_O; -- S msb) & O (lsb) -> D;/SP+1 
			when    RST_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & BLS_R & EXT_O; -- S->B; SP +1
			when    RST_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & PLD_P & NOP_A & SUP_R & EXT_O; -- S->P; SP+1
			when    RST_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SYU_R & EXT_O; -- S->Y (lsb); SP+1 (two byte instruction)  
			when    RST_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SYM_R & EXT_O; -- S->Y (msb); SP+1 (two byte instruction)  
			when    RST_OP7 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SXU_R & EXT_O; -- S->X (lsb); SP+1 (two byte instruction)
			when    RST_OP8 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SXM_R & EXT_O; -- S->X (msb); SP+1 (two byte instruction)
			when    RST_OP9 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SAU_R & EXT_O; -- S->A (lsb); SP+1 (two byte instruction) 
			when   RST_OP10 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & ALM_R & EXT_O; -- S->A (msb); EI   (two byte instruction) 
			
			-- PLP
			when    PLP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & PLD_P & NOP_A & NOP_R & EXT_O; -- S->P; EI 

			-- PLD
			when    PLD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLD_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- S->O (lsb); SP+1
			when    PLD_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & D16_R & EXM_O; -- S msb) & O (lsb) -> D; 
		
			-- PLA
			when    PLA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLA_OP1 =>
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- S->A (lsb); EI 
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- SP->MP; SP+1
               end if;		
			when    PLA_OP2 =>
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- S->O (msb)
					end if;				 
			when    PLA_OP3 =>
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & ORD_O; -- O->A (msb/lsb)
					end if;				 

			-- PLX
			when    PLX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLX_OP1 =>
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- S->X (lsb); EI 
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- SP->MP; SP+1
               end if;		
			when    PLX_OP2 =>
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- S->O (msb)
					end if;				 
			when    PLX_OP3 =>
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & ORD_O; -- O->X (msb/lsb)
					end if;				 

			-- PLY
			when    PLY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLY_OP1 =>
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- S->Y (lsb); EI 
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- SP->MP; SP+1
               end if;		
			when    PLY_OP2 =>
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- S->O (msb)
					end if;				 
			when    PLY_OP3 =>
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & ORD_O; -- O->X (msb/lsb)
					end if;				 

			-- PLR (in native mode PLR pulls ALWAYS 16 bit registers)
			when    PLR_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP;     SP+1 (two byte instruction)
			when    PLR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SYU_R & EXT_O; -- S->Y (lsb); SP+1 (two byte instruction)  
			when    PLR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SYM_R & EXT_O; -- S->Y (msb); SP+1 (two byte instruction)  
			when    PLR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SXU_R & EXT_O; -- S->X (lsb); SP+1 (two byte instruction)
			when    PLR_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SXM_R & EXT_O; -- S->X (msb); SP+1 (two byte instruction)
			when    PLR_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SAU_R & EXT_O; -- S->A (lsb); SP+1 (two byte instruction) 
			when    PLR_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & ALM_R & EXT_O; -- S->A (msb); EI   (two byte instruction) 
			
			-- RTI
			when    RTI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- PC->MEM; MP=01XX (STACK)
			when    RTI_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & PLD_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; MEM->P; SP +1
			when    RTI_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; LSB->O;  
			when    RTI_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTI_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MSB->O;  
			when    RTI_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- MP->MEM; SP +1;
			when    RTI_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADSP & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; MEM->PBR;

			-- RTS
			when    RTS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTS_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; LSB->O;  
			when    RTS_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- MP->MEM; SP +1;
			when    RTS_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MEM->PC
			when    RTS_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC+1; PC->MEM; EI

			-- ASL (A)
			when    ASL_OP0 =>
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & SHL_A & ALL_R & ARD_O; -- A (lsb) SHIFT LEFT; EI
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & SHL_A & A16_R & ARD_O; -- A (msb/lsb) SHIFT LEFT; EI
		           end if;			  

			-- LSR (A)
			when    LSR_OP0 => 
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & SHR_A & ALL_R & ARD_O; -- A (lsb) SHIFT RIGHT; EI
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & SHR_A & A16_R & ARD_O; -- A (msb/lsb) SHIFT RIGHT; EI
					  end if;  
			
			-- ROL (A)
			when    ROL_OP0 => 
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & ROL_A & ALL_R & ARD_O; -- A (lsb) ROTATE LEFT; EI
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & ROL_A & A16_R & ARD_O; -- A (msb\lsb) ROTATE LEFT; EI
		           end if;			  

			-- ROR (A)
			when    ROR_OP0 => 
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & ROR_A & ALL_R & ARD_O; -- A (lsb) ROTATE RIGHT; EI
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & ROR_A & A16_R & ARD_O; -- A (msb\lsb) ROTATE RIGHT; EI
		           end if;			  

			-- EXT (A)
			when    EXT_OP0 =>
			        if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- NOP; EI        (two byte instruction)
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & EXT_A & A16_R & ARD_O; -- A (msb/lsb) SHIFT LEFT; EI (two byte instruction)
		           end if;			  

			-- NEG (A)
			when    NEG_OP0 => 
			        if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NEG_A & ALL_R & ARD_O; -- negates A (lsb); EI (two byte instruction) 
					  else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NEG_A & A16_R & ARD_O; -- negates A (msb\lsb); EI (two byte instruction)
		           end if;			  
					  
			-- XYX
			when    XYX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & XRD_O; -- X->O;          (two byte instruction)
	  		when    XYX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & X16_R & YRD_O; -- Y->X; 
			when    XYX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NOP_A & Y16_R & ORD_O; -- O->Y; EI

			-- XAX
			when    XAX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & XRD_O; -- X->O;          (two byte instruction)
			when    XAX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & X16_R & ARD_O; -- A->X; 
			when    XAX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NOP_A & A16_R & ORD_O; -- O->A; EI

			-- XAY
			when    XAY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & YRD_O; -- Y->O;          (two byte instruction)
			when    XAY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & Y16_R & ARD_O; -- A->Y; 
			when    XAY_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NOP_A & A16_R & ORD_O; -- O->A; EI

			-- TCS  
			when    TCS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & S16_R & ARD_O; -- C->S;

			-- TSC  
			when    TSC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & SRD_O; -- S->C;
			
			-- XCE
			when    XCE_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & XCE_P & NOP_A & NOP_R & EXT_O; -- E<>C; EI

		   -- WDM
			when    WDM_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDM_P & NOP_A & NOP_R & EXT_O; -- set two byte instruction bit

			-- PHK
			when    PHK_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & KRD_O; -- K->S; SP-1; EI 
			
			-- PHB
			when    PHB_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & BRD_O; -- B->S; SP-1; EI 

			-- PLB
			when    PLB_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLB_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & BLD_R & EXT_O; -- S->B; EI 

			-- RTL
			when    RTL_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTL_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; LSB->O;  
			when    RTL_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTL_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MSB->O;  
			when    RTL_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- MP->MEM; SP +1;
			when    RTL_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; MEM->PBR;
			when    RTL_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC+1; PC->MEM; EI

			-- XBA
			when    XBA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & ARM_O; -- swap A<->B; EI

			-- WAI
			when    WAI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & WAI_R & EXT_O; -- set WAI flipflop
			when    WAI_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI

			-- STP
			when    STP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & STP_R & EXT_O; -- set STP flipflop
			when    STP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
			
			------------------------------------
			--           IMMEDIATE            --
			------------------------------------
			-- LDA #xx/#xxxx
			when  IMLDA_OP0 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MEM->A (lsb); PC +1; EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O (lsb); PC +1; EI
               end if;					
			when  IMLDA_OP1 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
					             q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MEM->A (msb\lsb); PC +1; EI
               end if;					
			
			-- LDX #xx/#xxxx
			when  IMLDX_OP0 => 
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MEM->X (lsb); PC +1; EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O (lsb); PC +1; EI
					end if;				 
			when  IMLDX_OP1 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else					
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & X16_R & EXM_O; -- MEM->X (msb\lsb); PC +1; EI
					end if;				 
					

			-- LDY #yy/#xxxx
			when  IMLDY_OP0 => 
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MEM->Y (lsb); PC +1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O (lsb); PC +1; EI
               end if;					
			when  IMLDY_OP1 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & Y16_R & EXM_O; -- MEM->Y (msb\lsb); PC +1; EI
					end if;				 

			-- ADC #xx/#xxxx (immediate)
			when  IMADC_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; PC +1; EI (emulation mode)
					else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); PC +1;
					end if;				 
			when  IMADC_OP1 =>  
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
				   else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
				   end if;					 
					
					
			-- SBC #xx/#xxxx (immediate)
			when  IMSBC_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-EXT; PC +1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- A=A+EXT; PC +1;
               end if;					
			when  IMSBC_OP1 =>
		         if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- MEM->A (msb\lsb); PC +1; EI
               end if;					

			-- CMP #xx/#xxxx (immediate)
			when  IMCMP_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM; PC +1; EI
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;;
               end if;	
			when  IMCMP_OP1 =>
		         if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-(msb\lsb); PC +1; EI
               end if;					

			-- CPX #xx/#xxxx (immediate)
			when  IMCPX_OP0 => 
			      if x = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-MEM; PC +1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;
               end if;	
			when  IMCPX_OP1 =>
		         if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-(msb\lsb); PC +1; EI
               end if;					
					

			-- CPY #xx/#xxxx (immediate)
			when  IMCPY_OP0 =>
			      if x = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y-MEM; PC +1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;
               end if;	
			when  IMCPY_OP1 =>
		         if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- X-(msb\lsb); PC +1; EI
               end if;					

			-- AND #xx/#xxxx (immediate)
			when  IMAND_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A AND MEM -> A; PC +1;
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;
               end if;	
		   when 	IMAND_OP1 => 
		         if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A AND MEM ->A (msb\lsb) -> A; PC +1; EI
               end if;					

			-- ORA #xx/#xxxx (immediate)
			when  IMORA_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A AND MEM -> A; PC +1;
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;
               end if;	
		   when 	IMORA_OP1 => 
		         if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A OR MEM ->A (msb\lsb) -> A; PC +1; EI
               end if;					

			-- EOR #xx (immediate)
			when  IMEOR_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A XOR MEM -> A; PC +1;
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;
               end if;	
		   when 	IMEOR_OP1 => 
		         if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A XOR MEM ->A (msb\lsb) -> A; PC +1; EI
               end if;					

			-- BIT #xx/#xxxx (immediate)
			when  IMBIT_OP0 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & LDZ_P & BIT_A & NOP_R & ARD_O; -- A AND MEM -> A; PC +1;
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM (lsb)->O; PC +1;
               end if;	
		   when 	IMBIT_OP1 => 
		         if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A AND MEM ->A (msb\lsb) -> A; PC +1; EI
               end if;					

			-- SEP #xx (immediate)
			when  IMSEP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & SEP_P & NOP_A & NOP_R & EXT_O; -- P = P OR MEM; PC +1;

			-- REP #xx (immediate)
			when  IMREP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & REP_P & NOP_A & NOP_R & EXT_O; -- P = P AND NOT MEM; PC +1;
			
			------------------------------------
			--           ZERO PAGE            --
			------------------------------------
			-- LDA $xx (zero page)      
			when  ZPLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLDA_OP1 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					 
			when  ZPLDA_OP2 => 
               if m = '1' then			
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1; EI
               end if;					

			-- LDX $xx (zero page)      
			when  ZPLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLDX_OP1 =>  
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZPLDX_OP2 => 
               if x = '1' then			
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & EXM_O; -- MP->MEM; MEM->X; PC+1; EI
               end if;					

			-- LDY $xx (zero page)      
			when  ZPLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLDY_OP1 => 
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZPLDY_OP2 => 
               if x = '1' then			
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & EXM_O; -- MP->MEM; MEM->Y; PC+1; EI
               end if;					

			-- STA $xx (zero page)      
			when  ZPSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTA_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A (lsb) ->MEM; PC+1; MP+1;
					end if;
			when  ZPSTA_OP2 =>
		         if m = '1' then 	
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A (msb) ->MEM; EI
               end if;					

			-- STX $xx (zero page)      
			when  ZPSTX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTX_OP1 => 
			      if x = '1' then  
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X->MEM; PC+1; EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X (lsb) ->MEM; PC+1; MP+1
					end if;
			when  ZPSTX_OP2 =>
		         if x = '1' then 	
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRM_O; -- MP->MEM; X (msb) ->MEM; EI
               end if;					
					

			-- STY $xx (zero page)      
			when  ZPSTY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTY_OP1 => 
			      if x = '1' then 
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y (lsb) ->MEM; PC+1; MP+1
					end if;
			when  ZPSTY_OP2 =>
		         if x = '1' then 	
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRM_O; -- MP->MEM; X (msb) ->MEM; EI;
               end if;					
					

			-- STZ $xx (zero page)      
			when  ZPSTZ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTZ_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; PC+1; EI
		         else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0 (lsb) ->MEM; PC+1; MP+1
               end if;					
			when  ZPSTZ_OP2 =>
		         if m = '1' then 	
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0 (msb) ->MEM; EI;
               end if;					
					
			-- ADC $xx (zero page)
			when  ZPADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPADC_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZPADC_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;

			-- SBC $xx (zero page)
			when  ZPSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSBC_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ZPSBC_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A - MEM(msb)\O(lsb) => A (msb\lsb); EI
               end if;

			-- CMP $xx (zeropage)
			when  ZPCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPCMP_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM; EI
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPCMP_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- CPX $xx (zeropage)
			when  ZPCPX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPCPX_OP1 => 
			      if x = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-MEM; EI
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPCPX_OP2 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X - MEM(msb)\O(lsb); EI
               end if;

			-- CPY $xx (zeropage)
			when  ZPCPY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPCPY_OP1 => 
			      if x = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y-MEM; EI
			      else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPCPY_OP2 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y - MEM(msb)\O(lsb); EI
               end if;

			-- AND $xx (zeropage)
			when  ZPAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPAND_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM;  EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPAND_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A = A AND MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xx (zeropage)
			when  ZPORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPORA_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM;  EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPORA_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A = A OR MEM(msb)\O(lsb); EI
               end if;

			-- EOR $xx (zeropage)
			when  ZPEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPEOR_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM;  EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPEOR_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A = A XOR MEM(msb)\O(lsb); EI
               end if;

			-- BIT $xx (zero page)      
			when  ZPBIT_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPBIT_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A BIT MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZPBIT_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A BIT MEM(msb)\O(lsb); EI
               end if;

			-- ASL $xx (zero page)
			when  ZPASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPASL_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPASL_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O SHIFT LEFT;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZPASL_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & SHL_A & O16_R & ORD_O; -- O SHIFT LEFT; MP-1
               end if;					
			when  ZPASL_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZPASL_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;

			-- LSR $xx (zero page)
			when  ZPLSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLSR_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPLSR_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O SHIFT RIGHT
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZPLSR_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & SHR_A & O16_R & ORD_O; -- O SHIFT LEFT; MP-1
               end if;					
			when  ZPLSR_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZPLSR_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;
			
			-- ROL $xx (zero page)
			when  ZPROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPROL_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPROL_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O ROTATE LEFT;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZPROL_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & ROL_A & O16_R & ORD_O; -- O ROTATE LEFT; MP-1
               end if;					
			when  ZPROL_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZPROL_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;
			
			-- ROR $xx (zero page)
			when  ZPROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPROR_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPROR_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O ROTATE RIGHT
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZPROR_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & ROR_A & O16_R & ORD_O; -- O ROTATE RIGHT; MP-1
               end if;					
			when  ZPROR_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZPROR_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;
			
			-- INC $xx (zero page)
			when  ZPINC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPINC_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPINC_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZPINC_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLD_P & INC_A & O16_R & ORD_O; -- O = O +1; MP-1
               end if;					
			when  ZPINC_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZPINC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;
			
			-- DEC $xx (zero page)
			when  ZPDEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPDEC_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPDEC_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O = O -1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (msb);
               end if;					
			when  ZPDEC_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLD_P & DEC_A & O16_R & ORD_O; -- O = O -1; MP-1
               end if;					
			when  ZPDEC_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZPDEC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;
			
			-- TSB $xx (zero page)
			when  ZPTSB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPTSB_OP1 =>
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPTSB_OP2 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> Z
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (msb);
               end if;		
			when  ZPTSB_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & TSB_A & OLD_R & ARD_O; -- A OR O -> O;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & LDZ_P & AND_A & O16_R & ARD_O; -- A AND O -> Z;
               end if;					
			when  ZPTSB_OP4 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & NOP_P & TSB_A & O16_R & ARD_O; -- A OR O -> O; MP -1
               end if;					
			when  ZPTSB_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; 
               end if;					
			when  ZPTSB_OP6 => 
               if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
               end if;					

			-- TRB $xx (zero page)
			when  ZPTRB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPTRB_OP1 =>
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZPTRB_OP2 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> Z
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (msb);
               end if;		
			when  ZPTRB_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & TRB_A & OLD_R & ARD_O; -- A NAND O -> O;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & LDZ_P & AND_A & O16_R & ARD_O; -- A AND O -> Z;
               end if;					
			when  ZPTRB_OP4 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & NOP_P & TRB_A & O16_R & ARD_O; -- A NAND O -> O; MP -1
               end if;					
			when  ZPTRB_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; 
               end if;					
			when  ZPTRB_OP6 => 
               if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
               end if;					
			
			------------------------------------
			--          ZERO PAGE,X           --  
			------------------------------------
			-- LDA $xx,X (zero page indexed)
			when  ZXLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXLDA_OP1 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; MP+1
               end if;					 
			when  ZXLDA_OP2 => 
               if m = '1' then			
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; EI
               end if;					
					
			-- LDY $xx,X (zero page indexed)
			when  ZXLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXLDY_OP1 => 
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXLDY_OP2 => 
               if x = '1' then			
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
				   else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & EXM_O; -- MP->MEM; MEM->Y; PC+1; EI
               end if;					
					
			-- STA $xx,X (zero page indexed)
			when  ZXSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSTA_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP+1
               end if;					
			when  ZXSTA_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; EI
               end if;					
					
			-- STY $xx,X (zero page indexed)
			when  ZXSTY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSTY_OP1 => 
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y->MEM; MP +1
               end if;					
			when  ZXSTY_OP2 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRM_O; -- MP->MEM; Y->MEM; EI
               end if;					
					
			-- STZ $xx,X (zero page indexed)
			when  ZXSTZ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSTZ_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; MP+1
               end if;					
			when  ZXSTZ_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; EI
               end if;					
					
			-- ADC $xx,X (zero page indexed)
			when  ZXADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXADC_OP1 => 
			      if m = '1' then 
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXADC_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
			
			-- SBC $xx,X (zero page indexed)
			when  ZXSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSBC_OP1 => 
			      if m = '1' then 
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXSBC_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
					
			-- CMP $xx,X (zero page indexed)
			when  ZXCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXCMP_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXCMP_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;
					
			-- AND $xx,X (zero page indexed)
			when  ZXAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXAND_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM;  EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXAND_OP2 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A - AND O -> A (msb/lsb); EI
               end if;
					
			-- ORA $xx,X (zero page indexed)
			when  ZXORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXORA_OP1 => 
			      if m = '1' then 
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM;  EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXORA_OP2 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A - OR O -> A (msb/lsb); EI
               end if;

			-- EOR $xx,X (zero page indexed)
			when  ZXEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXEOR_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM;  EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;					
			when  ZXEOR_OP2 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A - XOR O -> A (msb/lsb); EI
               end if;

			-- ASL $xx,X (zero page indexed)
			when  ZXASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXASL_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZXASL_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O SHIFT LEFT;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZXASL_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & SHL_A & O16_R & ORD_O; -- O SHIFT LEFT; MP-1
               end if;					
			when  ZXASL_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZXASL_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;
			
			-- LSR $xx,X (zero page indexed)
			when  ZXLSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXLSR_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZXLSR_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O SHIFT RIGHT
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZXLSR_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & SHR_A & O16_R & ORD_O; -- O SHIFT LEFT; MP-1
               end if;					
			when  ZXLSR_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZXLSR_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;

			-- ROL $xx,X (zero page indexed)
			when  ZXROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXROL_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZXROL_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O ROTATE LEFT;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZXROL_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & ROL_A & O16_R & ORD_O; -- O ROTATE LEFT; MP-1
               end if;					
			when  ZXROL_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZXROL_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;

			-- ROR $xx,X (zero page indexed)
			when  ZXROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXROR_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZXROR_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O ROTATE RIGHT
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZXROR_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLC_P & ROR_A & O16_R & ORD_O; -- O ROTATE RIGHT; MP-1
               end if;					
			when  ZXROR_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZXROR_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;

			-- INC $xx,X (zero page indexed)
			when  ZXINC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXINC_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZXINC_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
               end if;					
			when  ZXINC_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLD_P & INC_A & O16_R & ORD_O; -- O = O +1; MP-1
               end if;					
			when  ZXINC_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZXINC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;

			-- DEC $xx,X (zero page indexed)
			when  ZXDEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXDEC_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; MP +1
               end if;					
			when  ZXDEC_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O = O -1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O (msb);
               end if;					
			when  ZXDEC_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & DEC_M & FLD_P & DEC_A & O16_R & ORD_O; -- O = O -1; MP-1
               end if;					
			when  ZXDEC_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O(lsb)->MEM; MP +1
					end if;				 
			when  ZXDEC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O(msb)->MEM; EI
					end if;

			-- BIT $xx,X (zero page indexed)
			when  ZXBIT_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXBIT_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A BIT MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1; EI
               end if;
			when  ZXBIT_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A BIT MEM(msb)\O(lsb); EI
               end if;

			
			------------------------------------
			--          ZERO PAGE,Y           --
			------------------------------------
			-- LDX $xx,Y (zero page indexed)
			when  ZYLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZYLDX_OP1 => 
			      if x = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP +1
               end if;	
			when  ZYLDX_OP2 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O
               end if;	
			when  ZYLDX_OP3 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & ORD_O; -- O->X
               end if;	

			-- STX $xx,Y (zero page indexed)
			when  ZYSTX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZYSTX_OP1 => 
			      if x = '1' then 
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADDI & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X->MEM; MP +1
               end if;					
			when  ZYSTX_OP2 => 
			      if x = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRM_O; -- MP->MEM; X->MEM; EI
               end if;					
					

			------------------------------------
			--           INDIRECT             --
			------------------------------------
			-- JMP ($xxxx) (indirect)
			when  INJMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  INJMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  INJMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
			when  INJMP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MEM->PC; O->PC; EI

			-- JML ($xxxx) (indirect)
			when  INJML_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  INJML_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  INJML_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
			when  INJML_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
			when  INJML_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; EXT->PBR; EI
			
			------------------------------------
			--          INDIRECT,Y            --
			------------------------------------
			-- LDA ($xx),Y (zeropage - indirect - indexed)
			when  IYLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYLDA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYLDA_OP3 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  IYLDA_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;					
					
			-- STA ($xx),Y (zeropage - indirect - indexed)
			when  IYSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYSTA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYSTA_OP3 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP +1
               end if;					
			when  IYSTA_OP5 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; EI
               end if;					

			-- ADC ($xx),Y (zeropage - indirect - indexed)
			when  IYADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYADC_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  IYADC_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- A=A+MEM (msb)/O (lsb); EI
					end if;				 

			-- SBC ($xx),Y (zeropage - indirect - indexed)
			when  IYSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYSBC_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  IYSBC_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
					end if;

			-- CMP ($xx),Y (zeropage - indirect - indexed)
			when  IYCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYCMP_OP3 => 
			      if m = '1' then 
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM;  A-MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  IYCMP_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
					end if;

			-- AND ($xx),Y (zeropage - indirect - indexed)
			when  IYAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYAND_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  IYAND_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM (msb)/O (lsb); EI
					end if;

			-- ORA ($xx),Y (zeropage - indirect - indexed)
			when  IYORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYORA_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  IYORA_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM (msb)/O (lsb); EI
					end if;

			-- EOR ($xx),Y (zeropage - indirect - indexed)
			when  IYEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYEOR_OP3 => 
			      if m = '1' then 
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  IYEOR_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM (msb)/O (lsb); EI
					end if;
								 

			------------------------------------
			--          INDIRECT,X            --
			------------------------------------
			-- LDA ($xx,X) (zero page - indexed - indirect)
			when  IXLDA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXLDA_OP3 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI=1
					else				 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  IXLDA_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;					
			
			-- STA ($xx,X) (zero page - indexed - indirect)
			when  IXSTA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXSTA_OP3 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- A->MEM; EI=1
					else
 			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP +1
               end if;					
			when  IXSTA_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; EI
               end if;					

			-- AND ($xx,X) (zero page - indexed - indirect)
			when  IXAND_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXAND_OP3 => 
			      if m = '1' then 
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- MP->MEM; A=A AND MEM; EI=1
					else				 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  IXAND_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM (msb)/O (lsb); EI
					end if;

			-- ORA ($xx,X) (zero page - indexed - indirect)
			when  IXORA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXORA_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- MP->MEM; A=A OR MEM; EI=1
					else				 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  IXORA_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM (msb)/O (lsb); EI
					end if;

			-- EOR ($xx,X) (zero page - indexed - indirect)
			when  IXEOR_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXEOR_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- MP->MEM; A=A XOR MEM; EI=1
					else				 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  IXEOR_OP4 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM (msb)/O (lsb); EI
					end if;

			-- ADC ($xx,X) (zero page - indexed - indirect)
			when  IXADC_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXADC_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A + MEM; EI=1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  IXADC_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- A=A+MEM (msb)/O (lsb); EI
               end if;					
			
			-- SBC ($xx,X) (zero page - indexed - indirect)
			when  IXSBC_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXSBC_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A XOR MEM; EI=1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  IXSBC_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
               end if;					

			-- CMP ($xx,X) (zero page - indexed - indirect)
			when  IXCMP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXCMP_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM; A-MEM; EI=1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  IXCMP_OP4 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM (msb)/O (lsb); EI
               end if;					

			-- JMP ($xxxx,X) (absolute indexed - indirect)
			when  IXJMP_OP0 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  IXJMP_OP1 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ALL_M & AUC_P & SWC_A & NOP_R & XRD_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  IXJMP_OP2 => q <= ORD_D &'1'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ICC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MP_MSB+CARRY, EI
			when  IXJMP_OP3 => q <= ORD_D &'1'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
			when  IXJMP_OP4 => q <= ORD_D &'1'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADMP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			-- JSR ($xxxx,X) (absolute indexed - indirect)
			when  IXJSR_OP0 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  IXJSR_OP1 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1; 
			when  IXJSR_OP2 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1; 
			when  IXJSR_OP3 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ALL_M & AUC_P & SWC_A & NOP_R & XRD_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  IXJSR_OP4 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  IXJSR_OP5 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			------------------------------------
			--           ABSOLUTE             --
			------------------------------------
			-- LDA $xxxx (absolute)
			when  ABLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLDA_OP2 => 
			      if m = '1' then 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A (lsb);
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;	
			when  ABLDA_OP3 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;	

			-- LDX $xxxx (absolute)
			when  ABLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLDX_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLDX_OP2 => 
			      if x = '1' then 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->A (lsb);
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;	
			when  ABLDX_OP3 => 
			      if x = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;	

			-- LDY $xxxx (absolute)
			when  ABLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLDY_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLDY_OP2 => 
			      if x = '1' then 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y (lsb);
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;	
			when  ABLDY_OP3 => 
			      if x = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & EXM_O; -- MP->MEM; MEM->Y; PC+1
               end if;	

			-- STA $xxxx (absolute)
			when  ABSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTA_OP2 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A (lsb) ->MEM;
               end if;
			when  ABSTA_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A (msb) ->MEM;
               end if;					
					
			-- STX $xxxx (absolute)
			when  ABSTX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTX_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTX_OP2 => 
			      if x = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X (lsb) ->MEM;
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X (lsb) ->MEM;
               end if;
			when  ABSTX_OP3 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRM_O; -- MP->MEM; X (msb) ->MEM;
               end if;					

			-- STY $xxxx (absolute)
			when  ABSTY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTY_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTY_OP2 => 
			      if x = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y (lsb) ->MEM;
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y (lsb) ->MEM;
               end if;
			when  ABSTY_OP3 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRM_O; -- MP->MEM; Y (msb) ->MEM;
               end if;					
			
			-- STZ $xxxx (absolute)
			when  ABSTZ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTZ_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTZ_OP2 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; PC+1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0 (lsb) ->MEM;
               end if;
			when  ABSTZ_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0 (msb) ->MEM;
               end if;					
			
			-- JMP $xxxx (absolute)
			when  ABJMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			-- JSR $xxxx (absolute)
			when  ABJSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJSR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1; 
			when  ABJSR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1; 
			when  ABJSR_OP3 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			-- BIT $xxxx (absolute)
			when  ABBIT_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABBIT_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABBIT_OP2 => 
			      if m = '1' then 
                            q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- MP->MEM; MEM->ALU; PC+1	            
		         else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;	
			when  ABBIT_OP3 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- MP->MEM; BIT  
               end if;	

			-- ADC $xxxx (absolute)
			when  ABADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABADC_OP2 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABADC_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
			
			-- SBC $xxxx (absolute)
			when  ABSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSBC_OP2 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABSBC_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A = A - MEM(msb)\O(lsb); EI
               end if;
			
			-- CMP $xxxx (absolute)
			when  ABCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABCMP_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABCMP_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- CPX $xxxx (absolute)
			when  ABCPX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABCPX_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABCPX_OP2 => 
			      if x = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABCPX_OP3 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-MEM(msb)\O(lsb); EI
               end if;

			-- CPY $xxxx (absolute)
			when  ABCPY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABCPY_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABCPY_OP2 => 
			      if x = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- X-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABCPY_OP3 => 
			      if x = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y-MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xxxx (absolute)
			when  ABORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABORA_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABORA_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM(msb)\O(lsb); EI
               end if;

			-- AND $xxxx (absolute)
			when  ABAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABAND_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABAND_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM(msb)\O(lsb); EI
               end if;
			
			-- EOR $xxxx (absolute)
			when  ABEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABEOR_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ABEOR_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM(msb)\O(lsb); EI
               end if;

			-- ASL $xxxx (absolute)
			when  ABASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABASL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABASL_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ABASL_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O (lsb) SHIFT LEFT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  ABASL_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & SHL_A & O16_R & ORD_O; -- O (msb\lsb) SHIFT LEFT -> O; MP-1
               end if;
			when  ABASL_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  ABASL_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
					
			-- LSR $xxxx (absolute)
			when  ABLSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLSR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLSR_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ABLSR_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O (lsb) SHIFT RIGHT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  ABLSR_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & SHR_A & O16_R & ORD_O; -- O (msb\lsb) SHIFT RIGHT -> O; MP-1
               end if;
			when  ABLSR_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  ABLSR_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
			
			-- ROL $xxxx (absolute)
			when  ABROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABROL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABROL_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ABROL_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O (lsb) ROTATE LEFT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  ABROL_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & ROL_A & O16_R & ORD_O; -- O (msb\lsb) ROTATE LEFT -> O; MP-1
               end if;
			when  ABROL_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  ABROL_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
			
			-- ROR $xxxx (absolute)
			when  ABROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABROR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABROR_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ABROR_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O (lsb) ROTATE RIGHT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  ABROR_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & ROR_A & O16_R & ORD_O; -- O (msb\lsb) ROTATE RIGHT -> O; MP-1
               end if;
			when  ABROR_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  ABROR_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
			
			-- INC $xxxx (absolute)
			when  ABINC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABINC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABINC_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ABINC_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O  = O +1 -> O (lsb)
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  ABINC_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLD_P & INC_A & O16_R & ORD_O; -- O = O +1 (msb\lsb) -> O; MP-1
               end if;
			when  ABINC_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  ABINC_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
			
			-- DEC $xxxx (absolute)
			when  ABDEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABDEC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABDEC_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  ABDEC_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O  = O -1 -> O (lsb)
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  ABDEC_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLD_P & DEC_A & O16_R & ORD_O; -- O = O -1 (msb\lsb) -> O; MP-1
               end if;
			when  ABDEC_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP+1
			when  ABDEC_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
			
			-- TSB $xxxx (absolute)
			when  ABTSB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABTSB_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABTSB_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
               end if;					
			when  ABTSB_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> O
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O;
					end if;				 
			when  ABTSB_OP4 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & TSB_A & OLD_R & ARD_O; -- A OR O => O
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & LDZ_P & AND_A & O16_R & ARD_O; -- A AND O -> O
               end if;					
			when  ABTSB_OP5 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & NOP_P & TSB_A & O16_R & ARD_O; -- A OR O => O; MP-1
				   end if;					 
			when  ABTSB_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP+1
			when  ABTSB_OP7 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- TRB $xxxx (absolute)
			when  ABTRB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABTRB_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABTRB_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
               end if;					
			when  ABTRB_OP3 => 
			      if m = '1' then 
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> O
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O;
					end if;				 
			when  ABTRB_OP4 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & TSB_A & OLD_R & ARD_O; -- A OR O => O
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & LDZ_P & AND_A & O16_R & ARD_O; -- A AND O -> O
               end if;					
			when  ABTRB_OP5 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & NOP_P & TRB_A & O16_R & ARD_O; -- A NAND O => O; MP-1
				   end if;					 
			when  ABTRB_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP+1
			when  ABTRB_OP7 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;
			
			------------------------------------
			--          ABSOLUTE,X            --
			------------------------------------
	      --                      DMUX: ALU operand #2 multiplexer
	      --                      |       AI: effective address is indexed (X or Y)
	      --                      |       |   VP: vector pull
	      --                      |       |   |   ML: memory lock            
	      --                      |       |   |   |   VPA: vali program address 
	      --                      |       |   |   |   |   VDA: valid data address 
	      --                      |       |   |   |   |   |   EI: end of microcode sequence (the hidden extra cycle it's always executed after this microinstruction) 
	      --                      |       |   |   |   |   |   |   W: read/write control
	      --                      |       |   |   |   |   |   |   |    CLI: clear interrupt request
	      --                      |       |   |   |   |   |   |   |    |    PD: PC/MP address output multiplexer select
	      --                      |       |   |   |   |   |   |   |    |    |      PCR: register PC (program counter)
	      --                      |       |   |   |   |   |   |   |    |    |      |        MPR: register MP (memory pointer)
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       P_OP: register P set/reset bit
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       ALUOP: ALU operation
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       REGOP: registers load/increment/decrement etc.
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       RSEL: registers output multiplexer select
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
		   --                      DMUX    AI  VP  ML VPA VDA  EI  W    CLI  PD     PCR      MPR     P_OP    ALUOP   REGOP   RSEL
			-- LDA $xxxx,X (absolute indexed)
			when  AXLDA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXLDA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXLDA_OP2 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  AXLDA_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; EI
               end if;					

			-- LDY $xxxx,X (absolute indexed)
			when  AXLDY_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXLDY_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXLDY_OP2 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y; EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  AXLDY_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & Y16_R & EXM_O; -- MP->MEM; MEM->Y; EI
               end if;					
			
			-- STA $xxxx,X (absolute indexed)
			when  AXSTA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXSTA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXSTA_OP2 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI
					else 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP+1
               end if;					
			when  AXSTA_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; MP+1
               end if;					
			
			-- STZ $xxxx,X (absolute indexed)
			when  AXSTZ_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXSTZ_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXSTZ_OP2 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; MP+1
               end if;					
			when  AXSTZ_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; EI
               end if;					

			-- ADC $xxxx,X (absolute indexed)
			when  AXADC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXADC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXADC_OP2 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXADC_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
					
			-- SBC $xxxx,X (absolute indexed)
			when  AXSBC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXSBC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXSBC_OP2 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXSBC_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A - MEM(msb)\O(lsb)=> A (msb\lsb); EI
               end if;
			
			-- CMP $xxxx,X (absolute indexed)
			when  AXCMP_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXCMP_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXCMP_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXCMP_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;
					
			-- INC $xxxx,X (absolute indexed)
			when  AXINC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXINC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXINC_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  AXINC_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1 -> O (lsb)
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  AXINC_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLD_P & INC_A & O16_R & ORD_O; -- O = O +1 (msb\lsb) -> O; MP-1
               end if;
			when  AXINC_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  AXINC_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- DEC $xxxx,X (absolute indexed)
			when  AXDEC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXDEC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXDEC_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  AXDEC_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O  = O -1 -> O (lsb)
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  AXDEC_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLD_P & DEC_A & O16_R & ORD_O; -- O = O -1 (msb\lsb) -> O; MP-1
               end if;
			when  AXDEC_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  AXDEC_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- ASL $xxxx,X (absolute indexed)
			when  AXASL_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXASL_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXASL_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  AXASL_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O (lsb) SHIFT LEFT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  AXASL_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & SHL_A & O16_R & ORD_O; -- O (msb\lsb) SHIFT LEFT -> O; MP-1
               end if;
			when  AXASL_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  AXASL_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- LSR $xxxx,X (absolute indexed)
			when  AXLSR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXLSR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXLSR_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  AXLSR_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O (lsb) SHIFT RIGHT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  AXLSR_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & SHR_A & O16_R & ORD_O; -- O (msb\lsb) SHIFT RIGHT -> O; MP-1
               end if;
			when  AXLSR_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  AXLSR_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- ROL $xxxx,X (absolute indexed)
			when  AXROL_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXROL_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXROL_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  AXROL_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O (lsb) ROTATE LEFT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  AXROL_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & ROL_A & O16_R & ORD_O; -- O (msb\lsb) ROTATE LEFT -> O; MP-1
               end if;
			when  AXROL_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  AXROL_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- ROR $xxxx,X (absolute indexed)
			when  AXROR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXROR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXROR_OP2 => 
			      if m = '1' then
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb);
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  AXROR_OP3 => 
			      if m = '1' then  
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O (lsb) ROTATE RIGHT;
					else
					             q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
               end if;					
			when  AXROR_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; PC+1
					else
			                   q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & DEC_M & FLC_P & ROR_A & O16_R & ORD_O; -- O (msb\lsb) ROTATE RIGHT -> O; MP-1
               end if;
			when  AXROR_OP5 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O (lsb) ->MEM; MP +1
			when  AXROR_OP6 => q <= NOP_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & OMD_O; -- MP->MEM; O (msb) ->MEM;

			-- AND $xxxx,X (absolute indexed)
			when  AXAND_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXAND_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXAND_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & NOP_R & ARD_O; -- A AND EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXAND_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & NOP_R & ARD_O; -- A AND MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xxxx,X (absolute indexed)
			when  AXORA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXORA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXORA_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & NOP_R & ARD_O; -- A OR EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXORA_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & NOP_R & ARD_O; -- A OR MEM(msb)\O(lsb); EI
               end if;

			-- EOR $xxxx,X (absolute indexed)
			when  AXEOR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXEOR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXEOR_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & NOP_R & ARD_O; -- A XOR EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXEOR_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & NOP_R & ARD_O; -- A XOR MEM(msb)\O(lsb); EI
               end if;

			-- BIT $xxxx,X (absolute indexed)
			when  AXBIT_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXBIT_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXBIT_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A BIT EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AXBIT_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A BIT MEM(msb)\O(lsb); EI
               end if;
			
			------------------------------------
			--          ABSOLUTE,Y            --
			------------------------------------
			-- LDA $xxxx,Y (absolute indexed)
			when  AYLDA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYLDA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYLDA_OP2 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  AYLDA_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; EI
               end if;					

			-- LDX $xxxx,Y (absolute indexed)
			when  AYLDX_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYLDX_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYLDX_OP2 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
					end if;				 
			when  AYLDX_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & EXM_O; -- MP->MEM; MEM->X; EI
               end if;					

			-- STA $xxxx,Y (absolute indexed)
			when  AYSTA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYSTA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYSTA_OP2 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI
					else 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP+1
               end if;					
			when  AYSTA_OP3 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; MP+1
               end if;					

			-- ADC $xxxx,Y (absolute indexed)
			when  AYADC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYADC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYADC_OP2 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AYADC_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;

			-- SBC $xxxx,Y (absolute indexed)
			when  AYSBC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYSBC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYSBC_OP2 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AYSBC_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A - MEM(msb)\O(lsb)=> A (msb\lsb); EI
               end if;

			-- CMP $xxxx,Y (absolute indexed)
			when  AYCMP_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYCMP_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AYCMP_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AYCMP_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- AND $xxxx,Y (absolute indexed)
			when  AYAND_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYAND_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYAND_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & NOP_R & ARD_O; -- A AND EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AYAND_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & NOP_R & ARD_O; -- A AND MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xxxx,Y (absolute indexed)
			when  AYORA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYORA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYORA_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & NOP_R & ARD_O; -- A OR EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AYORA_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & NOP_R & ARD_O; -- A OR MEM(msb)\O(lsb); EI
               end if;

			-- EOR $xxxx,Y (absolute indexed)
			when  AYEOR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYEOR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYEOR_OP2 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & NOP_R & ARD_O; -- A XOR EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AYEOR_OP3 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & NOP_R & ARD_O; -- A XOR MEM(msb)\O(lsb); EI
               end if;
		
			
			--------------------------------------
			--          ABSOLUTE LONG           --
			--------------------------------------
			-- JML $xxxxxx (absolute long)
			when  ABJML_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJML_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ABJML_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; EXT->PBR; EI
	
			-- JSL $xxxxxx (absolute long)
			when  ABJSL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJSL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ABJSL_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & KRD_O; -- PBR->S; SP-1; 
			when  ABJSL_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1; 
			when  ABJSL_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1; 
			when  ABJSL_OP5 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; EXT->PBR; EI
	
			------------------------------------
			--            RELATIVE            --
			------------------------------------
			-- BRA xx
			when    BRA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;
			
			-- BEQ xx
			when    BEQ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BNE xx
			when    BNE_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BCC xx
			when    BCC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BCS xx
			when    BCS_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BVC xx
			when    BVC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BVS xx
			when    BVS_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BPL xx
			when    BPL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BMI xx
			when    BMI_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-----------------------------------------
			--            RELATIVE LONG            --
			-----------------------------------------
			-- BRL xxxx
			when    BRL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb offset);
			when    BRL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRL_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset

         -------------------------------
         --           STACK           --
         -------------------------------
         -- PEA xxxx
         when    PEA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
         when    PEA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; PC+1
			when    PEA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & OMD_O; -- O (msb) ->S; SP-1;
			when    PEA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ORD_O; -- O (lsb) ->S; SP-1;

         -- PEI xx
			when    PEI_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when    PEI_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when    PEI_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when    PEI_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & OMD_O; -- O (msb) ->S; SP-1;
			when    PEI_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ORD_O; -- O (lsb) ->S; SP-1;

         -- PER xxxx
			when    PER_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb offset);
			when    PER_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (msb offset)
			when    PER_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & SWC_A & O16_R & PCR_O; -- O = O + PC
			when    PER_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & OMD_O; -- O (msb) ->S; SP-1;
			when    PER_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ORD_O; -- O (lsb) ->S; SP-1;

			----------------------------------
			--          DIRECT,Y            --
			----------------------------------
			-- LDA [$xx],Y (zeropage - direct long - indexed)
			when  DYLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYLDA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYLDA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYLDA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MPR MSB
			when  DYLDA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYLDA_OP5 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  DYLDA_OP6 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;					
 
 			-- STA [$xx],Y (zeropage - indirect long - indexed)
			when  DYSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYSTA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYSTA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYSTA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYSTA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYSTA_OP5 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP +1
               end if;					
			when  DYSTA_OP6 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; EI
               end if;					

			-- ADC [$xx],Y (zeropage - indirect long - indexed)
			when  DYADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYADC_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYADC_OP5 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  DYADC_OP6 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- A=A+MEM (msb)/O (lsb); EI
					end if;				 

			-- SBC [$xx],Y (zeropage - indirect long - indexed)
			when  DYSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYSBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYSBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYSBC_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYSBC_OP5 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  DYSBC_OP6 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
					end if;

			-- CMP [$xx],Y (zeropage - indirect long - indexed)
			when  DYCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYCMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYCMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYCMP_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYCMP_OP5 => 
			      if m = '1' then 
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM;  A-MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DYCMP_OP6 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
					end if;

			-- AND [$xx],Y (zeropage - indirect long - indexed)
			when  DYAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYAND_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYAND_OP5 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DYAND_OP6 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM (msb)/O (lsb); EI
					end if;

			-- ORA [$xx],Y (zeropage - indirect long - indexed)
			when  DYORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYORA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYORA_OP5 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DYORA_OP6 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM (msb)/O (lsb); EI
					end if;

			-- EOR [$xx],Y (zeropage - indirect long - indexed)
			when  DYEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYEOR_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYEOR_OP5 => 
			      if m = '1' then 
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DYEOR_OP6 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM (msb)/O (lsb); EI
					end if;

			--------------------------------
			--          DIRECT            --
			--------------------------------
			-- LDA [$xx] (zeropage - direct long)
			when  DILDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DILDA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DILDA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DILDA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DILDA_OP4 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  DILDA_OP5 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;					
 
 			-- STA [$xx] (zeropage - indirect long)
			when  DISTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DISTA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DISTA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DISTA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DISTA_OP4 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; MP +1
               end if;					
			when  DISTA_OP5 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A->MEM; EI
               end if;					

			-- ADC [$xx] (zeropage - indirect long)
			when  DIADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIADC_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  DIADC_OP5 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- A=A+MEM (msb)/O (lsb); EI
					end if;				 

			-- SBC [$xx] (zeropage - indirect long)
			when  DISBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DISBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DISBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DISBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DISBC_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  DISBC_OP5 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
					end if;

			-- CMP [$xx] (zeropage - indirect long)
			when  DICMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DICMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DICMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DICMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DICMP_OP4 => 
			      if m = '1' then 
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM;  A-MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DICMP_OP5 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A=A-MEM (msb)/O (lsb); EI
					end if;

			-- AND [$xx] (zeropage - indirect long)
			when  DIAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIAND_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DIAND_OP5 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM (msb)/O (lsb); EI
					end if;

			-- ORA [$xx] (zeropage - indirect long)
			when  DIORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIORA_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DIORA_OP5 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM (msb)/O (lsb); EI
					end if;

			-- EOR [$xx] (zeropage - indirect long)
			when  DIEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIEOR_OP4 => 
			      if m = '1' then 
			                   q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;
			when  DIEOR_OP5 => 
			      if m = '1' then 
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else				 
			                   q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM (msb)/O (lsb); EI
					end if;
	
			----------------------------------------
			--           ABSOLUTE LONG            --
			----------------------------------------
			-- LDA $xxxxxx (absolute long)
			when  ALLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALLDA_OP3 => 
			      if m = '1' then 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A (lsb);
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;	
			when  ALLDA_OP4 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;	

			-- STA $xxxxxx (absolute long)
			when  ALSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALSTA_OP3 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A (lsb) ->MEM;
               end if;
			when  ALSTA_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A (msb) ->MEM;
               end if;					

			-- ADC $xxxxxx (absolute long)
			when  ALADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALADC_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ALADC_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
			
			-- SBC $xxxxxx (absolute long)
			when  ALSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALSBC_OP3 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ALSBC_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A = A - MEM(msb)\O(lsb); EI
               end if;
			
			-- CMP $xxxxxx (absolute long)
			when  ALCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALCMP_OP3 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ALCMP_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xxxxxx (absolute long)
			when  ALORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALORA_OP3 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ALORA_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM(msb)\O(lsb); EI
               end if;

			-- AND $xxxxxx (absolute long)
			when  ALAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALAND_OP3 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ALAND_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM(msb)\O(lsb); EI
               end if;
			
			-- EOR $xxxxxx (absolute long)
			when  ALEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALEOR_OP3 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  ALEOR_OP4 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM(msb)\O(lsb); EI
               end if;

			------------------------------------------
			--           ABSOLUTE LONG,X            --
			------------------------------------------
			-- LDA $xxxxxx,X (absolute long indexed X)
			when  AILDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AILDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AILDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AILDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AILDA_OP4 => 
			      if m = '1' then 
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A (lsb);
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;	
			when  AILDA_OP5 => 
			      if m = '1' then 
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
	            else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;	

			-- STA $xxxxxx,X (absolute long indexed X)
			when  AISTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AISTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AISTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AISTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AISTA_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A (lsb) ->MEM;
               end if;
			when  AISTA_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A (msb) ->MEM;
               end if;					
					
      	-- ADC $xxxxxx,X (absolute long indexed X)
			when  AIADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIADC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIADC_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AIADC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
			
			-- SBC $xxxxxx,X (absolute long indexed X)
			when  AISBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AISBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AISBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AISBC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AISBC_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AISBC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A = A - MEM(msb)\O(lsb); EI
               end if;
			
			-- CMP $xxxxxx,X (absolute long indexed X)
			when  AICMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AICMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AICMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AICMP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AICMP_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AICMP_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xxxxxx,X (absolute long indexed X)
			when  AIORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIORA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIORA_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AIORA_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM(msb)\O(lsb); EI
               end if;

			-- AND $xxxxxx,X (absolute long indexed X)
			when  AIAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIAND_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIAND_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AIAND_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM(msb)\O(lsb); EI
               end if;
			
			-- EOR $xxxxxx,X (absolute long indexed X)
			when  AIEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIEOR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIEOR_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  AIEOR_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM(msb)\O(lsb); EI
               end if;
					
			----------------------------------------
			--          STACK RELATIVE            --
			----------------------------------------
			-- LDA $xx,S (S + offset)
			when  SRLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRLDA_OP1 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  SRLDA_OP2 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;					

			-- STA $xx,S (S + offset)
			when  SRSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRSTA_OP1 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A (lsb) ->MEM;
               end if;
			when  SRSTA_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A (msb) ->MEM;
               end if;					

			-- ADC $xx,S (S + offset)
			when  SRADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRADC_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SRADC_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;
			
			-- SBC $xx,S (S + offset)
			when  SRSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRSBC_OP1 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SRSBC_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A = A - MEM(msb)\O(lsb); EI
               end if;
			
			-- CMP $xx,S (S + offset)
			when  SRCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRCMP_OP1 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SRCMP_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- ORA $xx,S (S + offset)
			when  SRORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRORA_OP1 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SRORA_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM(msb)\O(lsb); EI
               end if;

			-- AND $xx,S (S + offset)
			when  SRAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRAND_OP1 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SRAND_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM(msb)\O(lsb); EI
               end if;
			
			-- EOR $xx,S (S + offset)
			when  SREOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SREOR_OP1 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SREOR_OP2 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM(msb)\O(lsb); EI
               end if;
					
			-------------------------------------------------
			--          STACK RELATIVE INDEXED Y           --
			-------------------------------------------------
			-- LDA ($xx,S),Y
			when  SYLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYLDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYLDA_OP4 => 
			      if m = '1' then
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb); MP+1
               end if;					
			when  SYLDA_OP5 => 
			      if m = '1' then
			                   q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & EXM_O; -- MP->MEM; MEM->A; PC+1
               end if;					

			-- STA ($xx,S),Y
			when  SYSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYSTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYSTA_OP4 => 
			      if m = '1' then
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1
					else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A (lsb) ->MEM;
               end if;
			when  SYSTA_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
                            q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARM_O; -- MP->MEM; A (msb) ->MEM;
               end if;					

			-- ADC ($xx,S),Y
			when  SYADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYADC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYADC_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SYADC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & A16_R & ARD_O; -- MEM(msb)\O(lsb) + A => A (msb\lsb); PC +1; EI
               end if;

			-- SBC ($xx,S),Y
			when  SYSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYSBC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYSBC_OP4 => 
			      if m = '1' then
			                   q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SYSBC_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & A16_R & ARD_O; -- A = A - MEM(msb)\O(lsb); EI
               end if;

			-- CMP ($xx,S),Y
			when  SYCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYCMP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYCMP_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SYCMP_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A - MEM(msb)\O(lsb); EI
               end if;

			-- ORA ($xx,S),Y
			when  SYORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYORA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYORA_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SYORA_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & A16_R & ARD_O; -- A=A OR MEM(msb)\O(lsb); EI
               end if;

			-- AND ($xx,S),Y
			when  SYAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYAND_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYAND_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SYAND_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & A16_R & ARD_O; -- A=A AND MEM(msb)\O(lsb); EI
               end if;

			-- EOR ($xx,S),Y
			when  SYEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYEOR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYEOR_OP4 => 
			      if m = '1' then
					             q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI
               else
			                   q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM=>O (lsb); MP +1;
               end if;					
			when  SYEOR_OP5 => 
			      if m = '1' then
                            q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
               else
					             q <= EXM_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & A16_R & ARD_O; -- A=A XOR MEM(msb)\O(lsb); EI
               end if;
					
			------------------------------------
			--          MOVE BLOCK            --
			------------------------------------
         when  MBMVN_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (source)
			when  MBMVN_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADXR & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; read byte
         when  MBMVN_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (destination)
         when  MBMVN_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADYR & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O->MEM; write byte
         when  MBMVN_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MVN_R & EXT_O; -- X +1; Y +1; A -1;
         when  MBMVN_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & DE3_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- check for A = $FFFF 

         when  MBMVP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (source)
			when  MBMVP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADXR & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; read byte
         when  MBMVP_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (destination)
         when  MBMVP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADYR & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O->MEM; write byte
         when  MBMVP_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MVP_R & EXT_O; -- X -1; Y -1; A -1;
         when  MBMVP_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & DE3_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- check for A = $FFFF 
			
			----------------------------------
			--          MULTIPLY            --
			----------------------------------
			when    MPU_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MUI_R & EXT_O; -- load A/B & X on multiplier
			when    MPU_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MUS_R & EXT_O; -- start multiplication (unsigned)
			when    MPU_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & MUF_P & NOP_A & MUL_R & EXT_O; -- load result on A/B and X
			when    MPU_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- EI

			when    MPS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MUI_R & EXT_O; -- load A/B & X on multiplier
			when    MPS_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MSS_R & EXT_O; -- start multiplication (signed)
			when    MPS_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & MSF_P & NOP_A & MUL_R & EXT_O; -- load result on A/B and X
			when    MPS_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- EI
			
			when    others  => q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI

		end case;
	  else	 
		 -----------------------------------
		 --        EMULATION MODE         --
		 -----------------------------------
	    --                        DMUX: ALU operand #2 multiplexer
	    --                        |       AI: effective address is indexed (X or Y)
	    --                        |       |   VP: vector pull
	    --                        |       |   |   ML: memory lock            
	    --                        |       |   |   |   VPA: vali program address 
	    --                        |       |   |   |   |   VDA: valid data address 
	    --                        |       |   |   |   |   |   EI: end of microcode sequence (the hidden extra cycle it's always executed after this microinstruction) 
	    --                        |       |   |   |   |   |   |   W: read/write control
	    --                        |       |   |   |   |   |   |   |    CLI: clear interrupt request
	    --                        |       |   |   |   |   |   |   |    |    PD: PC/MP address output multiplexer select
	    --                        |       |   |   |   |   |   |   |    |    |      PCR: register PC (program counter)
	    --                        |       |   |   |   |   |   |   |    |    |      |        MPR: register MP (memory pointer)
	    --                        |       |   |   |   |   |   |   |    |    |      |        |       P_OP: register P set/reset bit
	    --                        |       |   |   |   |   |   |   |    |    |      |        |       |       ALUOP: ALU operation
	    --                        |       |   |   |   |   |   |   |    |    |      |        |       |       |       REGOP: registers load/increment/decrement etc.
	    --                        |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       RSEL: registers output multiplexer select
	    --                        |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
	    --                        |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
		 case a is              -- DMUX    AI  VP  ML VPA VDA  EI  W    CLI  PD     PCR      MPR     P_OP    ALUOP   REGOP   RSEL
			------------------------------------
			--            IMPLIED             --
			------------------------------------
			-- BRK
			when    BRK_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & IN2_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- if no interrupt request then PC=PC+2 
			when    BRK_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1 
			when    BRK_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1 
			when    BRK_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & VEC_M & SID_P & NOP_A & SDW_R & PRD_O; -- VEC->MP; SEI; CLD; 1->B (stack); P->S;
			when    BRK_OP4 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'0'& RDE &'1'& ADMP & LSB_PC & INC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCL; MP+1; interrupt ack; VP
			when    BRK_OP5 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'1'& RDE &'1'& ADMP & MSB_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCH; EI; VP 

			-- COP
			when    COP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & IN2_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC=PC+2 
			when    COP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1 
			when    COP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRL &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1 
			when    COP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & VEC_M & SID_P & NOP_A & SDW_R & PRD_O; -- VEC->MP; SEI; CLD; 1->B (stack); P->S;
			when    COP_OP4 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'0'& RDE &'1'& ADMP & LSB_PC & INC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCL; MP+1; interrupt ack; VP
			when    COP_OP5 => q <= ORD_D &'0'&'1'&'0'&'0'&'1'&'1'& RDE &'1'& ADMP & MSB_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->PCH; EI; VP 
			
			-- NOP
		   when    NOP_OP0 => q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
			
			-- CLC
			when    CLC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLC_P & NOP_A & NOP_R & EXT_O; -- 0->C; EI

			-- SEC
			when    SEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & SEC_P & NOP_A & NOP_R & EXT_O; -- 1->C; EI

			-- CLI
			when    CLI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLI_P & NOP_A & NOP_R & EXT_O; -- 0->I; EI

			-- SEI
			when    SEI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & SEI_P & NOP_A & NOP_R & EXT_O; -- 1->I; EI

			-- CLV
			when    CLV_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLV_P & NOP_A & NOP_R & EXT_O; -- 0->V; EI
			
			-- CLD
			when    CLD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & CLD_P & NOP_A & NOP_R & EXT_O; -- 0->D; EI

			-- SED
			when    SED_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & SED_P & NOP_A & NOP_R & EXT_O; -- 1->D; EI

			-- TAX
			when    TAX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & ARD_O; -- A->X; EI

			-- TXA
			when    TXA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & XRD_O; -- X->A; EI

			-- TAY
			when    TAY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & ARD_O; -- A->Y; EI

			-- TYA
			when    TYA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & YRD_O; -- Y->A; EI

			-- TXY
			when    TXY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & XRD_O; -- X->Y; EI

			-- TYX
			when    TYX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & YRD_O; -- Y->X; EI

			-- TCD
			when    TCD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & D16_R & ARD_O; -- C->D; EI

			-- TDC
			when    TDC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & DRD_O; -- D->C; EI

			-- TXS
			when    TXS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & S16_R & XRD_O; -- X->S; EI

			-- TSX
			when    TSX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & X16_R & SRD_O; -- S->X; EI

			-- INC A
			when    INC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & ALL_R & ARD_O; -- A+1; EI

			-- DEC A
			when    DEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & ALL_R & ARD_O; -- A-1; EI
			
			-- INX
			when    INX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & XLL_R & XRD_O; -- X+1; EI

			-- DEX
			when    DEX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & XLL_R & XRD_O; -- X-1; EI
			
			-- INY
			when    INY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & INC_A & YLL_R & YRD_O; -- Y+1; EI

			-- DEY
			when    DEY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & DEC_A & YLL_R & YRD_O; -- Y-1; EI

			-- PHP
			when    PHP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PRD_O; -- P->S; SP-1; EI 

			-- PHD
			when    PHD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & DRM_O; -- D (msb) ->S; SP-1;
			when    PHD_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & DRD_O; -- D (lsb) ->S; SP-1; EI 
		
			-- PHA
			when    PHA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A->S; SP-1; EI 

			-- PHX
			when    PHX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X->S; SP-1; EI 

			-- PHY
			when    PHY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRD_O; -- X->S; SP-1; EI 

			-- PHR (in emulation mode PHR pushes ALWAYS XY 8 bit registers and A as 16 bit register)
			when    PHR_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARM_O; -- A(msb)->S; SP-1;  (two byte instruction) 
			when    PHR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A(lsb)->S; SP-1;  (two byte instruction) 
			when    PHR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X->S; SP-1;       (two byte instruction)
			when    PHR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & SDW_R & YRD_O; -- Y->S; SP-1; EI    (two byte instruction)

			-- PLP
			when    PLP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & PLD_P & NOP_A & NOP_R & EXT_O; -- S->P; EI 

			-- SAV (in emulation mode SAV pushes ALWAYS XY 8 bit registers and A as 16 bit register)
			when    SAV_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARM_O; -- A(msb)->S; SP-1;  (two byte instruction) 
			when    SAV_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ARD_O; -- A(lsb)->S; SP-1;  (two byte instruction) 
			when    SAV_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & XRD_O; -- X->S; SP-1;     (two byte instruction)
			when    SAV_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & YRD_O; -- Y->S; SP-1;     (two byte instruction)
			when    SAV_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & BRD_O; -- B->S; SP-1;          (two byte instruction)
			when    SAV_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & DRM_O; -- D (msb) ->S; SP-1;   (two byte instruction)
			when    SAV_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & SDW_R & DRD_O; -- D (lsb) ->S; SP-1;   (two byte instruction)

			-- RST (in emulation mode RST pulls ALWAYS AXY 8 bit registers)
			when    RST_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP;     SP+1 (two byte instruction)
			when    RST_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- S->O (lsb); SP+1
			when    RST_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & DLS_R & EXM_O; -- S msb) & O (lsb) -> D;/SP+1 
			when    RST_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & BLS_R & EXT_O; -- S->B; SP +1
			when    RST_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SYU_R & EXT_O; -- S->Y;            (two byte instruction)  
			when    RST_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SXU_R & EXT_O; -- S->X;            (two byte instruction)
			when    RST_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SAU_R & EXT_O; -- S->A (lsb); SP+1 (two byte instruction) 
			when    RST_OP7 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & ALM_R & EXT_O; -- S->A (msb); EI   (two byte instruction) 
			
			-- PLD
			when    PLD_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLD_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OSU_R & EXT_O; -- S->O (lsb); SP+1
			when    PLD_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & D16_R & EXM_O; -- S msb) & O (lsb) -> D; 
			
			-- PLA
			when    PLA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- S->A; EI 

			-- PLX
			when    PLX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- S->X; EI 

			-- PLY
			when    PLY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- S->Y; EI 

			-- PLR (in emulation mode PLR pulls ALWAYS XY 8 bit registers and A as 16 bit register)
			when    PLR_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1     (two byte instruction)
			when    PLR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SYU_R & EXT_O; -- S->Y;            (two byte instruction)  
			when    PLR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SXU_R & EXT_O; -- S->X;            (two byte instruction)
			when    PLR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SAU_R & EXT_O; -- S->A (lsb); SP+1 (two byte instruction) 
			when    PLR_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & WDC_P & NOP_A & ALM_R & EXT_O; -- S->A (msb); EI   (two byte instruction) 
			
			-- RTI
			when    RTI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- PC->MEM; MP=01XX (STACK)
			when    RTI_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & PLD_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; MEM->P; SP +1
			when    RTI_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; LSB PC->O; SP +1; 
			when    RTI_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- MP->MEM; SP +1; 
			when    RTI_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; MSB->MP; EI

			-- RTS
			when    RTS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTS_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; LSB->O;  
			when    RTS_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- MP->MEM; SP +1;
			when    RTS_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MEM->PC
			when    RTS_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC+1; PC->MEM; EI

			-- ASL (A)
			when    ASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & SHL_A & ALL_R & ARD_O; -- A SHIFT LEFT; EI

			-- LSR (A)
			when    LSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & SHR_A & ALL_R & ARD_O; -- A SHIFT RIGHT; EI
			
			-- ROL (A)
			when    ROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & ROL_A & ALL_R & ARD_O; -- A ROTATE LEFT; EI

			-- ROR (A)
			when    ROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLC_P & ROR_A & ALL_R & ARD_O; -- A ROTATE RIGHT; EI

			-- EXT (A)
			when    EXT_OP0 => q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- NOP; EI        (two byte instruction)  
			
			-- NEG (A)
			when    NEG_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NEG_A & ALL_R & ARD_O; -- negates A (lsb); EI (two byte instruction)
			
			-- XYX
			when    XYX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & XRD_O; -- X->O;          (two byte instruction)
	  		when    XYX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & XLL_R & YRD_O; -- Y->X; 
			when    XYX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NOP_A & YLL_R & ORD_O; -- O->Y; EI

			-- XAX
			when    XAX_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & XRD_O; -- X->O;          (two byte instruction)
			when    XAX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & XLL_R & ARD_O; -- A->X; 
			when    XAX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NOP_A & ALL_R & ORD_O; -- O->A; EI

			-- XAY
			when    XAY_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & YRD_O; -- Y->O;          (two byte instruction)
			when    XAY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & YLL_R & ARD_O; -- A->Y; 
			when    XAY_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLW_P & NOP_A & ALL_R & ORD_O; -- O->A; EI

			-- TCS  
			when    TCS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & S16_R & ARD_O; -- C->S;

			-- TSC  
			when    TSC_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & SRD_O; -- S->C;
			
			-- XCE
			when    XCE_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & XCE_P & NOP_A & NOP_R & EXT_O; -- E-<>C; EI

		   -- WDM
			when    WDM_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDM_P & NOP_A & NOP_R & EXT_O; -- set two byte instruction bit

			-- PHK
			when    PHK_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & KRD_O; -- K->S; SP-1; EI 
			
			-- PHB
			when    PHB_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & BRD_O; -- B->S; SP-1; EI 

			-- PLB
			when    PLB_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MP; SP+1 
			when    PLB_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADSP & NOP_PC & NOP_M & FLD_P & NOP_A & BLD_R & EXT_O; -- S->B; EI 

			-- RTL
			when    RTL_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTL_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; LSB->O;  
			when    RTL_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- SP->MEM; SP +1
			when    RTL_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MSB->O;  
			when    RTL_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SUP_R & EXT_O; -- MP->MEM; SP +1;
			when    RTL_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADSP & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; MEM->PBR;
			when    RTL_OP6 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC+1; PC->MEM; EI

			-- XBA
			when    XBA_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLD_P & NOP_A & A16_R & ARM_O; -- swap A<->B; EI

			-- WAI
			when    WAI_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & WAI_R & EXT_O; -- set WAI flipflop
			when    WAI_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI

			-- STP
			when    STP_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & STP_R & EXT_O; -- set STP flipflop
			when    STP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
			
			------------------------------------
			--           IMMEDIATE            --
			------------------------------------
			-- LDA #xx
			when  IMLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MEM->A; PC +1; EI

			-- LDX #xx
			when  IMLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MEM->X; PC +1; EI

			-- LDY #yy
			when  IMLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MEM->Y; PC +1; EI

			-- ADC #xx (immediate)
			when  IMADC_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; PC +1; EI
			when  IMADC_OP1 => q <= BCD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAA_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); PC +1; EI

			-- SBC #xx (immediate)
			when  IMSBC_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-EXT; PC +1; EI
			when  IMSBC_OP1 => q <= BCD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAS_A & ALL_R & ARD_O; -- A=A-BCD ADJ (DAA); PC +1; EI

			-- CMP #xx (immediate)
			when  IMCMP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM; PC +1; EI

			-- CPX #xx (immediate)
			when  IMCPX_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-MEM; PC +1; EI

			-- CPY #xx (immediate)
			when  IMCPY_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y-MEM; PC +1; EI

			-- AND #xx (immediate)
			when  IMAND_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A AND MEM -> A; PC +1;

			-- ORA #xx (immediate)
			when  IMORA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A OR MEM -> A; PC +1;

			-- EOR #xx (immediate)
			when  IMEOR_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A XOR MEM -> A; PC +1;

			-- BIT #xx (immediate)
			when  IMBIT_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & LDZ_P & BIT_A & NOP_R & ARD_O; -- A AND MEM; PC +1;

			-- SEP #xx (immediate)
			when  IMSEP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & SEP_P &  OR_A & ALL_R & ARD_O; -- P = P OR MEM; PC +1;

			-- REP #xx (immediate)
			when  IMREP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & INC_PC & NOP_M & REP_P &  OR_A & ALL_R & ARD_O; -- P = P AND NOT MEM; PC +1;
			
			------------------------------------
			--           ZERO PAGE            --
			------------------------------------
			-- LDA $xx (zero page)      
			when  ZPLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; PC+1; EI

			-- LDX $xx (zero page)      
			when  ZPLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLDX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; PC+1; EI

			-- LDY $xx (zero page)      
			when  ZPLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLDY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y; PC+1; EI

			-- STA $xx (zero page)      
			when  ZPSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1; EI

			-- STX $xx (zero page)      
			when  ZPSTX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X->MEM; PC+1; EI

			-- STY $xx (zero page)      
			when  ZPSTY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y->MEM; PC+1; EI

			-- STZ $xx (zero page)      
			when  ZPSTZ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSTZ_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; PC+1; EI

			-- ADC $xx (zero page)
			when  ZPADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+MEM; EI
			when  ZPADC_OP2 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAA_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); PC +1; EI

			-- SBC $xx (zero page)
			when  ZPSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-MEM; EI
			when  ZPSBC_OP2 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAS_A & ALL_R & ARD_O; -- A=A-BCD ADJ (DAS); PC +1; EI

			-- CMP $xx (zeropage)
			when  ZPCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM; EI

			-- CPX $xx (zeropage)
			when  ZPCPX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPCPX_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-MEM; EI

			-- CPY $xx (zeropage)
			when  ZPCPY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPCPY_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y-MEM; EI

			-- AND $xx (zeropage)
			when  ZPAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM;  EI

			-- ORA $xx (zeropage)
			when  ZPORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM;  EI

			-- EOR $xx (zeropage)
			when  ZPEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM;  EI

			-- BIT $xx (zero page)      
			when  ZPBIT_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPBIT_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & INC_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- MP->MEM; MEM->ALU; PC+1; EI

			-- ASL $xx (zero page)
			when  ZPASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPASL_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPASL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O SHIFT LEFT;
			when  ZPASL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- LSR $xx (zero page)
			when  ZPLSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPLSR_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPLSR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O SHIFT RIGHT;
			when  ZPLSR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- ROL $xx (zero page)
			when  ZPROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPROL_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPROL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O ROTATE LEFT;
			when  ZPROL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- ROR $xx (zero page)
			when  ZPROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPROR_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPROR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O ROTATE RIGHT;
			when  ZPROR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- INC $xx (zero page)
			when  ZPINC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPINC_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPINC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1     
			when  ZPINC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- DEC $xx (zero page)
			when  ZPDEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPDEC_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPDEC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O = O -1    
			when  ZPDEC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- TSB $xx (zero page)
			when  ZPTSB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPTSB_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPTSB_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> Z
			when  ZPTSB_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & TSB_A & OLD_R & ARD_O; -- A OR O -> O
			when  ZPTSB_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI

			-- TRB $xx (zero page)
			when  ZPTRB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  ZPTRB_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1; EI
			when  ZPTRB_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> Z
			when  ZPTRB_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & TRB_A & OLD_R & ARD_O; -- A NAND O -> O
			when  ZPTRB_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1; EI
			
			------------------------------------
			--          ZERO PAGE,X           --  
			------------------------------------
			-- LDA $xx,X (zero page indexed)
			when  ZXLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI

			-- LDY $xx,X (zero page indexed)
			when  ZXLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXLDY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y; EI

			-- STA $xx,X (zero page indexed)
			when  ZXSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI

			-- STY $xx,X (zero page indexed)
			when  ZXSTY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSTY_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y->MEM; EI

			-- STZ $xx,X (zero page indexed)
			when  ZXSTZ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSTZ_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; X->MEM; EI

			-- ADC $xx,X (zero page indexed)
			when  ZXADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+MEM; EI
			when  ZXADC_OP2 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAA_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); EI

			-- SBC $xx,X (zero page indexed)
			when  ZXSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-MEM; EI
			when  ZXSBC_OP2 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAS_A & ALL_R & ARD_O; -- A=A-BCD ADJ (DAS); EI

			-- CMP $xx,X (zero page indexed)
			when  ZXCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-MEM; EI

			-- AND $xx,X (zero page indexed)
			when  ZXAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM;  EI

			-- ORA $xx,X (zero page indexed)
			when  ZXORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM;  EI

			-- EOR $xx,X (zero page indexed)
			when  ZXEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM;  EI

			-- ASL $xx,X (zero page indexed)
			when  ZXASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXASL_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; 
			when  ZXASL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O SHIFT LEFT;
			when  ZXASL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- LSR $xx,X (zero page indexed)
			when  ZXLSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXLSR_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
			when  ZXLSR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O SHIFT RIGHT;
			when  ZXLSR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- ROL $xx,X (zero page indexed)
			when  ZXROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXROL_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
			when  ZXROL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O ROTATE LEFT;
			when  ZXROL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- ROR $xx,X (zero page indexed)
			when  ZXROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXROR_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
			when  ZXROR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O ROTATE RIGHT;
			when  ZXROR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- INC $xx,X (zero page indexed)
			when  ZXINC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXINC_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
			when  ZXINC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1 
			when  ZXINC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- DEC $xx,X (zero page indexed)
			when  ZXDEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXDEC_OP1 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O;
			when  ZXDEC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O = O -1 
			when  ZXDEC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- BIT $xx,X (zero page indexed)
			when  ZXBIT_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZXBIT_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- A = A AND MEM;  EI
			
			------------------------------------
			--          ZERO PAGE,Y           --
			------------------------------------
			-- LDX $xx,Y (zero page indexed)
			when  ZYLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZYLDX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADDI & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; EI

			-- STX $xx,Y (zero page indexed)
			when  ZYSTX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & DOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+=D+O+X; PC+1;
			when  ZYSTX_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADDI & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X->MEM; EI

			------------------------------------
			--           INDIRECT             --
			------------------------------------
			-- JMP ($xxxx) (indirect)
			when  INJMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  INJMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  INJMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
			when  INJMP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MEM->PC; O->PC; EI

			-- JML ($xxxx) (indirect)
			when  INJML_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  INJML_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  INJML_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
			when  INJML_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MP->MEM; MEM->O; MP+1
			when  INJML_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; EXT->PBR; EI
			
			------------------------------------
			--          INDIRECT,Y            --
			------------------------------------
			-- LDA ($xx),Y (zeropage - indirect - indexed)
			when  IYLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYLDA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYLDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI

			-- STA ($xx),Y (zeropage - indirect - indexed)
			when  IYSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYSTA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYSTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI

			-- ADC ($xx),Y (zeropage - indirect - indexed)
			when  IYADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT

			-- SBC ($xx),Y (zeropage - indirect - indexed)
			when  IYSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYSBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT

			-- CMP ($xx),Y (zeropage - indirect - indexed)
			when  IYCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYCMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM;  A-MEM; EI

			-- AND ($xx),Y (zeropage - indirect - indexed)
			when  IYAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM; EI

			-- ORA ($xx),Y (zeropage - indirect - indexed)
			when  IYORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM; EI

			-- EOR ($xx),Y (zeropage - indirect - indexed)
			when  IYEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  IYEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  IYEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ABY_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O+Y->MP
			when  IYEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM; EI

			------------------------------------
			--          INDIRECT,X            --
			------------------------------------
			-- LDA ($xx,X) (zero page - indexed - indirect)
			when  IXLDA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB;
			when  IXLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXLDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI=1

			-- STA ($xx,X) (zero page - indexed - indirect)
			when  IXSTA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB;
			when  IXSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXSTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- A->MEM; EI=1

			-- AND ($xx,X) (zero page - indexed - indirect)
			when  IXAND_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB;
			when  IXAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- MP->MEM; A=A AND MEM; EI=1

			-- ORA ($xx,X) (zero page - indexed - indirect)
			when  IXORA_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB;
			when  IXORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- MP->MEM; A=A OR MEM; EI=1

			-- EOR ($xx,X) (zero page - indexed - indirect)
			when  IXEOR_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB;
			when  IXEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- MP->MEM; A=A XOR MEM; EI=1

			-- ADC ($xx,X) (zero page - indexed - indirect)
			when  IXADC_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB;
			when  IXADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A XOR MEM; EI=1
			when  IXADC_OP4 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAA_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); PC +1; EI

			-- SBC ($xx,X) (zero page - indexed - indirect)
			when  IXSBC_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXSBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A XOR MEM; EI=1
			when  IXSBC_OP4 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAS_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); PC +1; EI

			-- CMP ($xx,X) (zero page - indexed - indirect)
			when  IXCMP_OP0 => q <= EXT_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ZPL_M & NOP_P & SWC_A & NOP_R & XRD_O; -- ZP+X->MP; PC+1
			when  IXCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- O<=LSB; MP+=1
			when  IXCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ALL_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP<=MSB & LSB (O)
			when  IXCMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM; A=A XOR MEM; EI=1

			-- JMP ($xxxx,X) (absolute indexed - indirect)
			when  IXJMP_OP0 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  IXJMP_OP1 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ALL_M & AUC_P & SWC_A & NOP_R & XRD_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  IXJMP_OP2 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ICC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MEM->A; MP_MSB+CARRY, EI
			when  IXJMP_OP3 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  IXJMP_OP4 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			-- JSR ($xxxx,X) (absolute indexed - indirect)
			when  IXJSR_OP0 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  IXJSR_OP1 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1; 
			when  IXJSR_OP2 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1; 
			when  IXJSR_OP3 => q <= ORD_D &'1'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ALL_M & AUC_P & SWC_A & NOP_R & XRD_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  IXJSR_OP4 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  IXJSR_OP5 => q <= ORD_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			------------------------------------
			--           ABSOLUTE             --
			------------------------------------
			-- LDA $xxxx (absolute)
			when  ABLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; PC+1

			-- LDX $xxxx (absolute)
			when  ABLDX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLDX_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLDX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; PC+1

			-- LDY $xxxx (absolute)
			when  ABLDY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLDY_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLDY_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->Y; PC+1

			-- STA $xxxx (absolute)
			when  ABSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1

			-- STX $xxxx (absolute)
			when  ABSTX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTX_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & XRD_O; -- MP->MEM; X->MEM; PC+1

			-- STY $xxxx (absolute)
			when  ABSTY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTY_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTY_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & YRD_O; -- MP->MEM; Y->MEM; PC+1

			-- STZ $xxxx (absolute)
			when  ABSTZ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSTZ_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSTZ_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; PC+1
			
			-- JMP $xxxx (absolute)
			when  ABJMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			-- JSR $xxxx (absolute)
			when  ABJSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJSR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1; 
			when  ABJSR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1; 
			when  ABJSR_OP3 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LOD_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->PC; O->PC; EI

			-- BIT $xxxx (absolute)
			when  ABBIT_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABBIT_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABBIT_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- MP->MEM; MEM->ALU; PC+1

			-- ADC $xxxx (absolute)
			when  ABADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
			when  ABADC_OP3 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAA_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); PC +1; EI

			-- SBC $xxxx (absolute)
			when  ABSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABSBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A-EXT; EI
			when  ABSBC_OP3 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAS_A & ALL_R & ARD_O; -- A=A-BCD ADJ (DAA); PC +1; EI

			-- CMP $xxxx (absolute)
			when  ABCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABCMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI

			-- CPX $xxxx (absolute)
			when  ABCPX_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABCPX_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABCPX_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & XRD_O; -- X-EXT; EI

			-- CPY $xxxx (absolute)
			when  ABCPY_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABCPY_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABCPY_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & YRD_O; -- Y-EXT; EI

			-- ORA $xxxx (absolute)
			when  ABORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI

			-- AND $xxxx (absolute)
			when  ABAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI

			-- EOR $xxxx (absolute)
			when  ABEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI

			-- ASL $xxxx (absolute)
			when  ABASL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABASL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABASL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABASL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O SHIFT LEFT;
			when  ABASL_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- LSR $xxxx (absolute)
			when  ABLSR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABLSR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABLSR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABLSR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O SHIFT RIGHT;
			when  ABLSR_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- ROL $xxxx (absolute)
			when  ABROL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABROL_OP1 => q <= ORD_D &'0'&'0'&'1'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABROL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABROL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O ROTATE LEFT;
			when  ABROL_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- ROR $xxxx (absolute)
			when  ABROR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABROR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABROR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABROR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O ROTATE RIGHT;
			when  ABROR_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- INC $xxxx (absolute)
			when  ABINC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABINC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABINC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABINC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1
			when  ABINC_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- DEC $xxxx (absolute)
			when  ABDEC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABDEC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABDEC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABDEC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O = O -1
			when  ABDEC_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- TSB $xxxx (absolute)
			when  ABTSB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABTSB_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABTSB_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABTSB_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> Z
			when  ABTSB_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & TSB_A & OLD_R & ARD_O; -- A OR O => O
			when  ABTSB_OP5 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1

			-- TRB $xxxx (absolute)
			when  ABTRB_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & LSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- LSB->MP; PC+1
			when  ABTRB_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MSB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MSB->MP; PC+1
			when  ABTRB_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; PC+1
			when  ABTRB_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & LDZ_P & AND_A & NOP_R & ARD_O; -- A AND O -> Z
			when  ABTRB_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & TRB_A & OLD_R & ARD_O; -- A NAND O => O
			when  ABTRB_OP5 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; PC+1
			
			------------------------------------
			--          ABSOLUTE,X            --
			------------------------------------
	      --                      DMUX: ALU operand #2 multiplexer
	      --                      |       AI: effective address is indexed (X or Y)
	      --                      |       |   VP: vector pull
	      --                      |       |   |   ML: memory lock            
	      --                      |       |   |   |   VPA: vali program address 
	      --                      |       |   |   |   |   VDA: valid data address 
	      --                      |       |   |   |   |   |   EI: end of microcode sequence (the hidden extra cycle it's always executed after this microinstruction) 
	      --                      |       |   |   |   |   |   |   W: read/write control
	      --                      |       |   |   |   |   |   |   |    CLI: clear interrupt request
	      --                      |       |   |   |   |   |   |   |    |    PD: PC/MP address output multiplexer select
	      --                      |       |   |   |   |   |   |   |    |    |      PCR: register PC (program counter)
	      --                      |       |   |   |   |   |   |   |    |    |      |        MPR: register MP (memory pointer)
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       P_OP: register P set/reset bit
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       ALUOP: ALU operation
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       REGOP: registers load/increment/decrement etc.
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       RSEL: registers output multiplexer select
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
	      --                      |       |   |   |   |   |   |   |    |    |      |        |       |       |       |       |
		   --                      DMUX    AI  VP  ML VPA VDA  EI  W    CLI  PD     PCR      MPR     P_OP    ALUOP   REGOP   RSEL
			-- LDA $xxxx,X (absolute indexed)
			when  AXLDA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXLDA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXLDA_OP2 => q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
			
			-- LDY $xxxx,X (absolute indexed)
			when  AXLDY_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXLDY_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXLDY_OP2 => q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & YLL_R & EXT_O; -- MP->MEM; MEM->A; EI
			
			-- STA $xxxx,X (absolute indexed)
			when  AXSTA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXSTA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXSTA_OP2 => q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI

			-- STZ $xxxx,X (absolute indexed)
			when  AXSTZ_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXSTZ_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXSTZ_OP2 => q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & Z00_O; -- MP->MEM; 0->MEM; EI

			-- ADC $xxxx,X (absolute indexed)
			when  AXADC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXADC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT

			-- SBC $xxxx,X (absolute indexed)
			when  AXSBC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXSBC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXSBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT; EI
			
			-- CMP $xxxx,X (absolute indexed)
			when  AXCMP_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXCMP_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXCMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM; A-MEM MP_MSB+CARRY, EI

			-- INC $xxxx,X (absolute indexed)
			when  AXINC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXINC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXINC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  AXINC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & INC_A & OLD_R & ORD_O; -- O = O +1     
			when  AXINC_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- DEC $xxxx,X (absolute indexed)
			when  AXDEC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXDEC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXDEC_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  AXDEC_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & DEC_A & OLD_R & ORD_O; -- O = O -1     
			when  AXDEC_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- ASL $xxxx,X (absolute indexed)
			when  AXASL_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXASL_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXASL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  AXASL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHL_A & OLD_R & ORD_O; -- O SHIFT LEFT 
			when  AXASL_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- LSR $xxxx,X (absolute indexed)
			when  AXLSR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXLSR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXLSR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  AXLSR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & SHR_A & OLD_R & ORD_O; -- O SHIFT RIGHT
			when  AXLSR_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- ROL $xxxx,X (absolute indexed)
			when  AXROL_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXROL_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXROL_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  AXROL_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROL_A & OLD_R & ORD_O; -- O ROTATE LEFT 
			when  AXROL_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- ROR $xxxx,X (absolute indexed)
			when  AXROR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXROR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXROR_OP2 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O; EI
			when  AXROR_OP3 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & ROR_A & OLD_R & ORD_O; -- O ROTATE RIGHT
			when  AXROR_OP4 => q <= ORD_D &'0'&'0'&'1'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- MP->MEM; O->MEM; EI

			-- AND $xxxx,X (absolute indexed)
			when  AXAND_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXAND_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- MP->MEM; EXT AND A; EI

			-- ORA $xxxx,X (absolute indexed)
			when  AXORA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXORA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- MP->MEM; EXT OR A; EI

			-- EOR $xxxx,X (absolute indexed)
			when  AXEOR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXEOR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- MP->MEM; EXT XOR A; EI

			-- BIT $xxxx,X (absolute indexed)
			when  AXBIT_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AXBIT_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+X->MP_LSB; PC+1;
			when  AXBIT_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & BIT_A & NOP_R & ARD_O; -- MP->MEM; EXT BIT A; EI
			
			------------------------------------
			--          ABSOLUTE,Y            --
			------------------------------------
			-- LDA $xxxx,X (absolute indexed)
			when  AYLDA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYLDA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYLDA_OP2 => q <= NOP_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI

			-- LDX $xxxx,Y (absolute indexed)
			when  AYLDX_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYLDX_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYLDX_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & ICC_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; MP_MSB+CARRY, EI
			when  AYLDX_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & XLL_R & EXT_O; -- MP->MEM; MEM->X; EI

			-- STA $xxxx,Y (absolute indexed)
			when  AYSTA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYSTA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ICC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; MP_MSB+CARRY, EI
			when  AYSTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI

			-- ADC $xxxx,Y (absolute indexed)
			when  AYADC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYADC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ICC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; A=A+EXT; MP_MSB+CARRY, EI
			when  AYADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT
			when  AYADC_OP4 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAA_A & ALL_R & ARD_O; -- A=A+BCD ADJ (DAA); PC +1; EI

			-- SBC $xxxx,Y (absolute indexed)
			when  AYSBC_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYSBC_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYSBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ICC_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP->MEM; A=A-EXT; MP_MSB+CARRY, EI
			when  AYSBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT
			when  AYSBC_OP4 => q <= BCD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & FLV_P & DAS_A & ALL_R & ARD_O; -- A=A-BCD ADJ (DAS); PC +1; EI

			-- CMP $xxxx,Y (absolute indexed)
			when  AYCMP_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYCMP_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYCMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & ICC_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM; A-MEM MP_MSB+CARRY, EI
			when  AYCMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM; A-MEM; EI

			-- AND $xxxx,Y (absolute indexed)
			when  AYAND_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYAND_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & ICC_M & FLD_P & AND_A & ALL_R & ARD_O; -- MP->MEM; EXT AND A; MP_MSB+CARRY, EI
			when  AYAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- MP->MEM; EXT AND A; EI

			-- ORA $xxxx,Y (absolute indexed)
			when  AYORA_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYORA_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & ICC_M & FLD_P &  OR_A & ALL_R & ARD_O; -- MP->MEM; EXT OR A; MP_MSB+CARRY, EI
			when  AYORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- MP->MEM; EXT OR A; EI

			-- EOR $xxxx,Y (absolute indexed)
			when  AYEOR_OP0 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
			when  AYEOR_OP1 => q <= NOP_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & ABY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->MP_MSB; MEM->O+Y->MP_LSB; PC+1;
			when  AYEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & ICC_M & FLD_P & XOR_A & ALL_R & ARD_O; -- MP->MEM; EXT XOR A; MP_MSB+CARRY, EI
			when  AYEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- MP->MEM; EXT XOR A; EI

			--------------------------------------
			--          ABSOLUTE LONG           --
			--------------------------------------
			-- JML $xxxxxx (absolute long)
			when  ABJML_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJML_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ABJML_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; EXT->PRB; EI

			-- JSL $xxxxxx (absolute long)
			when  ABJSL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ABJSL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ABJSL_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & KRD_O; -- PBR->S; SP-1; 
			when  ABJSL_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PHR_O; -- PCH->S; SP-1; 
			when  ABJSL_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & PLR_O; -- PCL->S; SP-1; 
			when  ABJSL_OP5 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & LML_PC & NOP_M & NOP_P & NOP_A & KLD_R & EXT_O; -- O->PC; EXT->PBR; EI
			
			------------------------------------
			--            RELATIVE            --
			------------------------------------
			-- BRA xx
			when    BRA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;
			
			-- BEQ xx
			when    BEQ_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BNE xx
			when    BNE_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BCC xx
			when    BCC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BCS xx
			when    BCS_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BVC xx
			when    BVC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BVS xx
			when    BVS_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BPL xx
			when    BPL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-- BMI xx
			when    BMI_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRA_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset;

			-----------------------------------------
			--            RELATIVE LONG            --
			-----------------------------------------
			-- BRL xxxx
			when    BRL_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb offset);
			when    BRL_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'1'& RDE &'0'& ADPC & BRL_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- PC +1 + offset

         -------------------------------
         --           STACK           --
         -------------------------------
         -- PEA xxxx
         when    PEA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; PC+1
         when    PEA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; PC+1
			when    PEA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & OMD_O; -- O (msb) ->S; SP-1;
			when    PEA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ORD_O; -- O (lsb) ->S; SP-1;
			
         -- PEI xx
			when    PEI_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when    PEI_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when    PEI_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when    PEI_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & OMD_O; -- O (msb) ->S; SP-1;
			when    PEI_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ORD_O; -- O (lsb) ->S; SP-1;

         -- PER xxxx
			when    PER_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MP->MEM; MEM->O (lsb offset);
			when    PER_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (msb offset)
			when    PER_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & SWC_A & O16_R & PCR_O; -- O = O + PC
			when    PER_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & OMD_O; -- O (msb) ->S; SP-1;
			when    PER_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADSP & NOP_PC & NOP_M & NOP_P & NOP_A & SDW_R & ORD_O; -- O (lsb) ->S; SP-1;

			----------------------------------
			--          DIRECT,Y            --
			----------------------------------
			-- LDA [$xx],Y (zeropage - direct long - indexed)
			when  DYLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYLDA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYLDA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYLDA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYLDA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYLDA_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
 
 			-- STA [$xx],Y (zeropage - indirect long - indexed)
			when  DYSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYSTA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYSTA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYSTA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYSTA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYSTA_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI

			-- ADC [$xx],Y (zeropage - indirect long - indexed)
			when  DYADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYADC_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYADC_OP5 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT

			-- SBC [$xx],Y (zeropage - indirect long - indexed)
			when  DYSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYSBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYSBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYSBC_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYSBC_OP5 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT

			-- CMP [$xx],Y (zeropage - indirect long - indexed)
			when  DYCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYCMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYCMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYCMP_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYCMP_OP5 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM;  A-MEM; EI

			-- AND [$xx],Y (zeropage - indirect long - indexed)
			when  DYAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYAND_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYAND_OP5 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM; EI

			-- ORA [$xx],Y (zeropage - indirect long - indexed)
			when  DYORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYORA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYORA_OP5 => q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM; EI

			-- EOR [$xx],Y (zeropage - indirect long - indexed)
			when  DYEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DYEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DYEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DYEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DYEOR_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & ADY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  DYEOR_OP5 => q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM; EI

			--------------------------------
			--          DIRECT            --
			--------------------------------
			-- LDA [$xx] (zeropage - direct long)
			when  DILDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DILDA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DILDA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DILDA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
  		   when  DILDA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI
 
 			-- STA [$xx] (zeropage - indirect long)
			when  DISTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DISTA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DISTA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DISTA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DISTA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; EI

			-- ADC [$xx] (zeropage - indirect long)
			when  DIADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIADC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIADC_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- MP->MEM; A=A+EXT

			-- SBC [$xx] (zeropage - indirect long)
			when  DISBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DISBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DISBC_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DISBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DISBC_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- MP->MEM; A=A-EXT

			-- CMP [$xx] (zeropage - indirect long)
			when  DICMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DICMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DICMP_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DICMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DICMP_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- MP->MEM;  A-MEM; EI

			-- AND [$xx] (zeropage - indirect long)
			when  DIAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIAND_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIAND_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A = A AND MEM; EI

			-- ORA [$xx] (zeropage - indirect long)
			when  DIORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIORA_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIORA_OP4 => q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A = A OR MEM; EI

			-- EOR [$xx] (zeropage - indirect long)
			when  DIEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & ZPL_M & NOP_P & NOP_A & NOP_R & EXT_O; -- ZP->MP; PC+1
			when  DIEOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & INC_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; (LSB POINTER)
			when  DIEOR_OP2 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MEM->O; (MSB POINTER)
			when  DIEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MEM->B
			when  DIEOR_OP4 => q <= EXT_D &'1'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A = A XOR MEM; EI

			----------------------------------------
			--           ABSOLUTE LONG            --
			----------------------------------------
			-- LDA $xxxxxx (absolute long)
			when  ALLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALLDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A

			-- STA $xxxxxx (absolute long)
			when  ALSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALSTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; 

			-- ADC $xxxxxx (absolute long)
			when  ALADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALADC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
			
			-- SBC $xxxxxx (absolute long)
			when  ALSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALSBC_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
			
			-- CMP $xxxxxx (absolute long)
			when  ALCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALCMP_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI

			-- ORA $xxxxxx (absolute long)
			when  ALORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALORA_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI

			-- AND $xxxxxx (absolute long)
			when  ALAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALAND_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
			
			-- EOR $xxxxxx (absolute long)
			when  ALEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  ALEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  ALEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  ALEOR_OP3 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI

			------------------------------------------
			--           ABSOLUTE LONG,X            --
			------------------------------------------
			-- LDA $xxxxxx,X (absolute long indexed X)
			when  AILDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AILDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AILDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AILDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AILDA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A (lsb);

			-- STA $xxxxxx,X (absolute long indexed X)
			when  AISTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AISTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AISTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AISTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AISTA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1
					
			-- ADC $xxxxxx,X (absolute long indexed X)
			when  AIADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIADC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIADC_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
			
			-- SBC $xxxxxx,X (absolute long indexed X)
			when  AISBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AISBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AISBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AISBC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AISBC_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
			
			-- CMP $xxxxxx,X (absolute long indexed X)
			when  AICMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AICMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AICMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AICMP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AICMP_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI

			-- ORA $xxxxxx,X (absolute long indexed X)
			when  AIORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIORA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIORA_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI

			-- AND $xxxxxx,X (absolute long indexed X)
			when  AIAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIAND_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIAND_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
			
			-- EOR $xxxxxx,X (absolute long indexed X)
			when  AIEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; PC+1
			when  AIEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O; PC+1
			when  AIEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & MHB_M & NOP_P & NOP_A & NOP_R & EXT_O; -- HIGH->MP; PC+1
			when  AIEOR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & ADX_M & NOP_P & NOP_A & NOP_R & EXT_O; -- O+Y->MP (24 bit)
			when  AIEOR_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI

			----------------------------------------
			--          STACK RELATIVE            --
			----------------------------------------
			-- LDA $xx,S (S + offset)
			when  SRLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI

			-- STA $xx,S (S + offset)
			when  SRSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1

			-- ADC $xx,S (S + offset)
			when  SRADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRADC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI
			
			-- SBC $xx,S (S + offset)
			when  SRSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRSBC_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI
			
			-- CMP $xx,S (S + offset)
			when  SRCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRCMP_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI

			-- ORA $xx,S (S + offset)
			when  SRORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRORA_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI

			-- AND $xx,S (S + offset)
			when  SRAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SRAND_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI
			
			-- EOR $xx,S (S + offset)
			when  SREOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SREOR_OP1 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI

			-------------------------------------------------
			--          STACK RELATIVE INDEXED Y           --
			-------------------------------------------------
			-- LDA ($xx,S),Y
			when  SYLDA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYLDA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYLDA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYLDA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYLDA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & NOP_A & ALL_R & EXT_O; -- MP->MEM; MEM->A; EI

			-- STA ($xx,S),Y
			when  SYSTA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYSTA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYSTA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYSTA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYSTA_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'1'& WRE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ARD_O; -- MP->MEM; A->MEM; PC+1

			-- ADC ($xx,S),Y
			when  SYADC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYADC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYADC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYADC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYADC_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUM_A & ALL_R & ARD_O; -- A=A+EXT; EI

			-- SBC ($xx,S),Y
			when  SYSBC_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYSBC_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYSBC_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYSBC_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYSBC_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLV_P & SUB_A & ALL_R & ARD_O; -- A=A+EXT; EI

			-- CMP ($xx,S),Y
			when  SYCMP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYCMP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYCMP_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYCMP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYCMP_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLC_P & CMP_A & NOP_R & ARD_O; -- A-EXT; EI

			-- ORA ($xx,S),Y
			when  SYORA_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYORA_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYORA_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYORA_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYORA_OP5 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P &  OR_A & ALL_R & ARD_O; -- A=A OR MEM; EI

			-- AND ($xx,S),Y
			when  SYAND_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYAND_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYAND_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYAND_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYAND_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & AND_A & ALL_R & ARD_O; -- A=A AND MEM; EI

			-- EOR ($xx,S),Y
			when  SYEOR_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & AOS_M & NOP_P & NOP_A & NOP_R & EXT_O; -- S+OFFSET->MP; PC+1
			when  SYEOR_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & INC_M & NOP_P & NOP_A & OLD_R & EXT_O; -- LSB->O; MP+1
			when  SYEOR_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADMP & NOP_PC & NOP_M & NOP_P & NOP_A & OMD_R & EXT_O; -- MSB->O;
			when  SYEOR_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADMP & NOP_PC & AOY_M & NOP_P & NOP_A & NOP_R & EXT_O; -- MP+O+Y
			when  SYEOR_OP4 => q <= EXT_D &'0'&'0'&'0'&'0'&'1'&'1'& RDE &'0'& ADMP & NOP_PC & NOP_M & FLD_P & XOR_A & ALL_R & ARD_O; -- A=A XOR MEM; EI

			------------------------------------
			--          MOVE BLOCK            --
			------------------------------------
         when  MBMVN_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (source)
			when  MBMVN_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADXR & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; read byte
         when  MBMVN_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (destination)
         when  MBMVN_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADYR & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O->MEM; write byte
         when  MBMVN_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MVN_R & EXT_O; -- X +1; Y +1; A -1;
         when  MBMVN_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & DE3_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- check for A = $FFFF 

         when  MBMVP_OP0 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (source)
			when  MBMVP_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& RDE &'0'& ADXR & NOP_PC & NOP_M & NOP_P & NOP_A & OLD_R & EXT_O; -- MEM->O; read byte
         when  MBMVP_OP2 => q <= ORD_D &'0'&'0'&'0'&'1'&'0'&'0'& RDE &'0'& ADPC & INC_PC & NOP_M & NOP_P & NOP_A & BLD_R & EXT_O; -- MEM->DBR (destination)
         when  MBMVP_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'1'&'0'& WRE &'0'& ADYR & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & ORD_O; -- O->MEM; write byte
         when  MBMVP_OP4 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MVP_R & EXT_O; -- X -1; Y -1; A -1;
         when  MBMVP_OP5 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & DE3_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- check for A = $FFFF 

			----------------------------------
			--          MULTIPLY            --
			----------------------------------
   		when    MPU_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MUI_R & EXT_O; -- load A/B & X on multiplier
			when    MPU_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MUS_R & EXT_O; -- start multiplication (unsigned)
			when    MPU_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & MUF_P & NOP_A & MUL_R & EXT_O; -- load result on A/B and X
			when    MPU_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- EI

			when    MPS_OP0 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MUI_R & EXT_O; -- load A/B & X on multiplier
			when    MPS_OP1 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & MSS_R & EXT_O; -- start multiplication (signed)
			when    MPS_OP2 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'0'& RDE &'0'& ADPC & NOP_PC & NOP_M & MSF_P & NOP_A & MUL_R & EXT_O; -- load result on A/B and X
			when    MPS_OP3 => q <= ORD_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & WDC_P & NOP_A & NOP_R & EXT_O; -- EI
			
			when    others  => q <= NOP_D &'0'&'0'&'0'&'0'&'0'&'1'& RDE &'0'& ADPC & NOP_PC & NOP_M & NOP_P & NOP_A & NOP_R & EXT_O; -- EI
		 end case;
	  end if;		 
  end process;
end comb;


